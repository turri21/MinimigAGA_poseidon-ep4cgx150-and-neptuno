// minimig version constants

localparam [7:0] BETA_FLAG  = 8'd1;  // BETA / RELEASE flag
localparam [7:0] MAJOR_VER  = 8'd20;  // major version number (Year)
localparam [7:0] MINOR_VER  = 8'd09;  // minor version number (Month)
localparam [7:0] MINION_VER = 8'd15;  // least version number (Day)

