library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"01",
     1 => x"da",
     2 => x"87",
     3 => x"04",
     4 => x"dd",
     5 => x"87",
     6 => x"0e",
     7 => x"58",
     8 => x"5e",
     9 => x"59",
    10 => x"5a",
    11 => x"0e",
    12 => x"27",
    13 => x"00",
    14 => x"00",
    15 => x"00",
    16 => x"2c",
    17 => x"0f",
    18 => x"26",
    19 => x"4a",
    20 => x"26",
    21 => x"49",
    22 => x"26",
    23 => x"48",
    24 => x"ff",
    25 => x"80",
    26 => x"26",
    27 => x"08",
    28 => x"4f",
    29 => x"27",
    30 => x"00",
    31 => x"00",
    32 => x"00",
    33 => x"2d",
    34 => x"4f",
    35 => x"27",
    36 => x"00",
    37 => x"00",
    38 => x"00",
    39 => x"29",
    40 => x"4f",
    41 => x"00",
    42 => x"fd",
    43 => x"87",
    44 => x"4f",
    45 => x"c1",
    46 => x"cc",
    47 => x"e4",
    48 => x"4e",
    49 => x"c9",
    50 => x"c0",
    51 => x"86",
    52 => x"c1",
    53 => x"cc",
    54 => x"e4",
    55 => x"49",
    56 => x"c1",
    57 => x"c3",
    58 => x"c0",
    59 => x"48",
    60 => x"89",
    61 => x"d0",
    62 => x"89",
    63 => x"03",
    64 => x"c0",
    65 => x"40",
    66 => x"40",
    67 => x"40",
    68 => x"40",
    69 => x"f6",
    70 => x"87",
    71 => x"d0",
    72 => x"81",
    73 => x"05",
    74 => x"c0",
    75 => x"50",
    76 => x"c1",
    77 => x"89",
    78 => x"05",
    79 => x"f9",
    80 => x"87",
    81 => x"c1",
    82 => x"c3",
    83 => x"c0",
    84 => x"4d",
    85 => x"c1",
    86 => x"c3",
    87 => x"c0",
    88 => x"4c",
    89 => x"74",
    90 => x"ad",
    91 => x"02",
    92 => x"c4",
    93 => x"87",
    94 => x"24",
    95 => x"0f",
    96 => x"f7",
    97 => x"87",
    98 => x"c1",
    99 => x"c4",
   100 => x"87",
   101 => x"c1",
   102 => x"c3",
   103 => x"c0",
   104 => x"4d",
   105 => x"c1",
   106 => x"c3",
   107 => x"c0",
   108 => x"4c",
   109 => x"74",
   110 => x"ad",
   111 => x"02",
   112 => x"c6",
   113 => x"87",
   114 => x"c4",
   115 => x"8c",
   116 => x"6c",
   117 => x"0f",
   118 => x"f5",
   119 => x"87",
   120 => x"00",
   121 => x"fd",
   122 => x"87",
   123 => x"1e",
   124 => x"73",
   125 => x"1e",
   126 => x"c2",
   127 => x"c0",
   128 => x"c0",
   129 => x"4b",
   130 => x"73",
   131 => x"0f",
   132 => x"c4",
   133 => x"87",
   134 => x"26",
   135 => x"4d",
   136 => x"26",
   137 => x"4c",
   138 => x"26",
   139 => x"4b",
   140 => x"26",
   141 => x"4f",
   142 => x"1e",
   143 => x"71",
   144 => x"4a",
   145 => x"c0",
   146 => x"f6",
   147 => x"e4",
   148 => x"c0",
   149 => x"c4",
   150 => x"49",
   151 => x"c0",
   152 => x"e0",
   153 => x"9f",
   154 => x"79",
   155 => x"c0",
   156 => x"e1",
   157 => x"9f",
   158 => x"79",
   159 => x"c0",
   160 => x"e0",
   161 => x"9f",
   162 => x"79",
   163 => x"c0",
   164 => x"e1",
   165 => x"9f",
   166 => x"79",
   167 => x"26",
   168 => x"4f",
   169 => x"1e",
   170 => x"73",
   171 => x"1e",
   172 => x"c4",
   173 => x"fe",
   174 => x"49",
   175 => x"c0",
   176 => x"f1",
   177 => x"c4",
   178 => x"87",
   179 => x"c0",
   180 => x"fc",
   181 => x"c0",
   182 => x"4b",
   183 => x"cf",
   184 => x"e2",
   185 => x"87",
   186 => x"70",
   187 => x"98",
   188 => x"02",
   189 => x"c0",
   190 => x"f4",
   191 => x"87",
   192 => x"c0",
   193 => x"ff",
   194 => x"f0",
   195 => x"4b",
   196 => x"c4",
   197 => x"e7",
   198 => x"49",
   199 => x"c0",
   200 => x"f0",
   201 => x"ec",
   202 => x"87",
   203 => x"d5",
   204 => x"ed",
   205 => x"87",
   206 => x"70",
   207 => x"98",
   208 => x"02",
   209 => x"da",
   210 => x"87",
   211 => x"c3",
   212 => x"f0",
   213 => x"4b",
   214 => x"c2",
   215 => x"c0",
   216 => x"c0",
   217 => x"1e",
   218 => x"c3",
   219 => x"ff",
   220 => x"49",
   221 => x"c0",
   222 => x"ed",
   223 => x"df",
   224 => x"87",
   225 => x"c4",
   226 => x"86",
   227 => x"70",
   228 => x"98",
   229 => x"02",
   230 => x"cc",
   231 => x"87",
   232 => x"fe",
   233 => x"d0",
   234 => x"87",
   235 => x"c7",
   236 => x"87",
   237 => x"c4",
   238 => x"cb",
   239 => x"49",
   240 => x"c0",
   241 => x"f0",
   242 => x"c3",
   243 => x"87",
   244 => x"73",
   245 => x"49",
   246 => x"fe",
   247 => x"d5",
   248 => x"87",
   249 => x"fe",
   250 => x"f0",
   251 => x"87",
   252 => x"fe",
   253 => x"cb",
   254 => x"87",
   255 => x"38",
   256 => x"33",
   257 => x"32",
   258 => x"4f",
   259 => x"53",
   260 => x"44",
   261 => x"41",
   262 => x"41",
   263 => x"42",
   264 => x"49",
   265 => x"4e",
   266 => x"00",
   267 => x"55",
   268 => x"6e",
   269 => x"61",
   270 => x"62",
   271 => x"6c",
   272 => x"65",
   273 => x"20",
   274 => x"74",
   275 => x"6f",
   276 => x"20",
   277 => x"6c",
   278 => x"6f",
   279 => x"63",
   280 => x"61",
   281 => x"74",
   282 => x"65",
   283 => x"20",
   284 => x"70",
   285 => x"61",
   286 => x"72",
   287 => x"74",
   288 => x"69",
   289 => x"74",
   290 => x"69",
   291 => x"6f",
   292 => x"6e",
   293 => x"0a",
   294 => x"00",
   295 => x"48",
   296 => x"75",
   297 => x"6e",
   298 => x"74",
   299 => x"69",
   300 => x"6e",
   301 => x"67",
   302 => x"20",
   303 => x"66",
   304 => x"6f",
   305 => x"72",
   306 => x"20",
   307 => x"70",
   308 => x"61",
   309 => x"72",
   310 => x"74",
   311 => x"69",
   312 => x"74",
   313 => x"69",
   314 => x"6f",
   315 => x"6e",
   316 => x"0a",
   317 => x"00",
   318 => x"49",
   319 => x"6e",
   320 => x"69",
   321 => x"74",
   322 => x"69",
   323 => x"61",
   324 => x"6c",
   325 => x"69",
   326 => x"7a",
   327 => x"69",
   328 => x"6e",
   329 => x"67",
   330 => x"20",
   331 => x"53",
   332 => x"44",
   333 => x"20",
   334 => x"63",
   335 => x"61",
   336 => x"72",
   337 => x"64",
   338 => x"0a",
   339 => x"00",
   340 => x"1e",
   341 => x"e4",
   342 => x"86",
   343 => x"c0",
   344 => x"f6",
   345 => x"e4",
   346 => x"c0",
   347 => x"c0",
   348 => x"4a",
   349 => x"c3",
   350 => x"ff",
   351 => x"97",
   352 => x"7a",
   353 => x"97",
   354 => x"6a",
   355 => x"48",
   356 => x"c4",
   357 => x"a6",
   358 => x"58",
   359 => x"6e",
   360 => x"49",
   361 => x"c3",
   362 => x"ff",
   363 => x"99",
   364 => x"97",
   365 => x"7a",
   366 => x"c8",
   367 => x"31",
   368 => x"97",
   369 => x"6a",
   370 => x"48",
   371 => x"c8",
   372 => x"a6",
   373 => x"58",
   374 => x"c4",
   375 => x"66",
   376 => x"48",
   377 => x"c3",
   378 => x"ff",
   379 => x"98",
   380 => x"cc",
   381 => x"a6",
   382 => x"58",
   383 => x"c8",
   384 => x"66",
   385 => x"b1",
   386 => x"c3",
   387 => x"ff",
   388 => x"97",
   389 => x"7a",
   390 => x"c8",
   391 => x"31",
   392 => x"97",
   393 => x"6a",
   394 => x"48",
   395 => x"d0",
   396 => x"a6",
   397 => x"58",
   398 => x"cc",
   399 => x"66",
   400 => x"48",
   401 => x"c3",
   402 => x"ff",
   403 => x"98",
   404 => x"d4",
   405 => x"a6",
   406 => x"58",
   407 => x"d0",
   408 => x"66",
   409 => x"b1",
   410 => x"c3",
   411 => x"ff",
   412 => x"97",
   413 => x"7a",
   414 => x"c8",
   415 => x"31",
   416 => x"12",
   417 => x"48",
   418 => x"d8",
   419 => x"a6",
   420 => x"58",
   421 => x"d4",
   422 => x"66",
   423 => x"48",
   424 => x"c3",
   425 => x"ff",
   426 => x"98",
   427 => x"dc",
   428 => x"a6",
   429 => x"58",
   430 => x"d8",
   431 => x"66",
   432 => x"b1",
   433 => x"71",
   434 => x"48",
   435 => x"e4",
   436 => x"8e",
   437 => x"26",
   438 => x"4f",
   439 => x"0e",
   440 => x"5e",
   441 => x"5b",
   442 => x"5c",
   443 => x"5d",
   444 => x"0e",
   445 => x"1e",
   446 => x"71",
   447 => x"4a",
   448 => x"c0",
   449 => x"f6",
   450 => x"e4",
   451 => x"c0",
   452 => x"c0",
   453 => x"4b",
   454 => x"72",
   455 => x"49",
   456 => x"c3",
   457 => x"ff",
   458 => x"99",
   459 => x"73",
   460 => x"09",
   461 => x"97",
   462 => x"79",
   463 => x"09",
   464 => x"c1",
   465 => x"c3",
   466 => x"c0",
   467 => x"bf",
   468 => x"05",
   469 => x"c8",
   470 => x"87",
   471 => x"d4",
   472 => x"66",
   473 => x"48",
   474 => x"c9",
   475 => x"30",
   476 => x"d8",
   477 => x"a6",
   478 => x"58",
   479 => x"d4",
   480 => x"66",
   481 => x"49",
   482 => x"d8",
   483 => x"29",
   484 => x"c3",
   485 => x"ff",
   486 => x"99",
   487 => x"73",
   488 => x"09",
   489 => x"97",
   490 => x"79",
   491 => x"09",
   492 => x"d4",
   493 => x"66",
   494 => x"49",
   495 => x"d0",
   496 => x"29",
   497 => x"c3",
   498 => x"ff",
   499 => x"99",
   500 => x"73",
   501 => x"09",
   502 => x"97",
   503 => x"79",
   504 => x"09",
   505 => x"d4",
   506 => x"66",
   507 => x"49",
   508 => x"c8",
   509 => x"29",
   510 => x"c3",
   511 => x"ff",
   512 => x"99",
   513 => x"73",
   514 => x"09",
   515 => x"97",
   516 => x"79",
   517 => x"09",
   518 => x"d4",
   519 => x"66",
   520 => x"49",
   521 => x"c3",
   522 => x"ff",
   523 => x"99",
   524 => x"73",
   525 => x"09",
   526 => x"97",
   527 => x"79",
   528 => x"09",
   529 => x"72",
   530 => x"49",
   531 => x"d0",
   532 => x"29",
   533 => x"c3",
   534 => x"ff",
   535 => x"99",
   536 => x"73",
   537 => x"09",
   538 => x"97",
   539 => x"79",
   540 => x"09",
   541 => x"97",
   542 => x"6b",
   543 => x"48",
   544 => x"c4",
   545 => x"a6",
   546 => x"58",
   547 => x"6e",
   548 => x"4c",
   549 => x"c3",
   550 => x"ff",
   551 => x"9c",
   552 => x"c9",
   553 => x"f0",
   554 => x"ff",
   555 => x"4d",
   556 => x"c3",
   557 => x"ff",
   558 => x"ac",
   559 => x"05",
   560 => x"da",
   561 => x"87",
   562 => x"c3",
   563 => x"ff",
   564 => x"97",
   565 => x"7b",
   566 => x"97",
   567 => x"6b",
   568 => x"48",
   569 => x"c4",
   570 => x"a6",
   571 => x"58",
   572 => x"6e",
   573 => x"4c",
   574 => x"c3",
   575 => x"ff",
   576 => x"9c",
   577 => x"c1",
   578 => x"8d",
   579 => x"02",
   580 => x"c6",
   581 => x"87",
   582 => x"c3",
   583 => x"ff",
   584 => x"ac",
   585 => x"02",
   586 => x"e6",
   587 => x"87",
   588 => x"74",
   589 => x"4a",
   590 => x"c4",
   591 => x"b7",
   592 => x"2a",
   593 => x"c0",
   594 => x"f0",
   595 => x"a2",
   596 => x"49",
   597 => x"c0",
   598 => x"ea",
   599 => x"d0",
   600 => x"87",
   601 => x"74",
   602 => x"4a",
   603 => x"cf",
   604 => x"9a",
   605 => x"c0",
   606 => x"f0",
   607 => x"a2",
   608 => x"49",
   609 => x"c0",
   610 => x"ea",
   611 => x"c4",
   612 => x"87",
   613 => x"74",
   614 => x"48",
   615 => x"26",
   616 => x"26",
   617 => x"4d",
   618 => x"26",
   619 => x"4c",
   620 => x"26",
   621 => x"4b",
   622 => x"26",
   623 => x"4f",
   624 => x"1e",
   625 => x"c0",
   626 => x"49",
   627 => x"c0",
   628 => x"f6",
   629 => x"e4",
   630 => x"c0",
   631 => x"c0",
   632 => x"48",
   633 => x"c3",
   634 => x"ff",
   635 => x"50",
   636 => x"c1",
   637 => x"81",
   638 => x"c3",
   639 => x"c8",
   640 => x"b7",
   641 => x"a9",
   642 => x"04",
   643 => x"ee",
   644 => x"87",
   645 => x"26",
   646 => x"4f",
   647 => x"0e",
   648 => x"5e",
   649 => x"5b",
   650 => x"5c",
   651 => x"0e",
   652 => x"c0",
   653 => x"f6",
   654 => x"e4",
   655 => x"c0",
   656 => x"c0",
   657 => x"4c",
   658 => x"ff",
   659 => x"db",
   660 => x"87",
   661 => x"c4",
   662 => x"f8",
   663 => x"df",
   664 => x"4b",
   665 => x"c0",
   666 => x"1e",
   667 => x"c0",
   668 => x"ff",
   669 => x"f0",
   670 => x"c1",
   671 => x"f7",
   672 => x"49",
   673 => x"fc",
   674 => x"d3",
   675 => x"87",
   676 => x"c4",
   677 => x"86",
   678 => x"c1",
   679 => x"a8",
   680 => x"05",
   681 => x"c0",
   682 => x"e6",
   683 => x"87",
   684 => x"c3",
   685 => x"ff",
   686 => x"97",
   687 => x"7c",
   688 => x"c1",
   689 => x"c0",
   690 => x"c0",
   691 => x"c0",
   692 => x"c0",
   693 => x"c0",
   694 => x"1e",
   695 => x"c0",
   696 => x"e1",
   697 => x"f0",
   698 => x"c1",
   699 => x"e9",
   700 => x"49",
   701 => x"fb",
   702 => x"f7",
   703 => x"87",
   704 => x"c4",
   705 => x"86",
   706 => x"70",
   707 => x"98",
   708 => x"05",
   709 => x"c8",
   710 => x"87",
   711 => x"c3",
   712 => x"ff",
   713 => x"97",
   714 => x"7c",
   715 => x"c1",
   716 => x"48",
   717 => x"cb",
   718 => x"87",
   719 => x"fe",
   720 => x"de",
   721 => x"87",
   722 => x"c1",
   723 => x"8b",
   724 => x"05",
   725 => x"ff",
   726 => x"c1",
   727 => x"87",
   728 => x"c0",
   729 => x"48",
   730 => x"fe",
   731 => x"cd",
   732 => x"87",
   733 => x"43",
   734 => x"4d",
   735 => x"44",
   736 => x"34",
   737 => x"31",
   738 => x"20",
   739 => x"25",
   740 => x"64",
   741 => x"0a",
   742 => x"00",
   743 => x"43",
   744 => x"4d",
   745 => x"44",
   746 => x"35",
   747 => x"35",
   748 => x"20",
   749 => x"25",
   750 => x"64",
   751 => x"0a",
   752 => x"00",
   753 => x"43",
   754 => x"4d",
   755 => x"44",
   756 => x"34",
   757 => x"31",
   758 => x"20",
   759 => x"25",
   760 => x"64",
   761 => x"0a",
   762 => x"00",
   763 => x"43",
   764 => x"4d",
   765 => x"44",
   766 => x"35",
   767 => x"35",
   768 => x"20",
   769 => x"25",
   770 => x"64",
   771 => x"0a",
   772 => x"00",
   773 => x"69",
   774 => x"6e",
   775 => x"69",
   776 => x"74",
   777 => x"20",
   778 => x"25",
   779 => x"64",
   780 => x"0a",
   781 => x"20",
   782 => x"20",
   783 => x"00",
   784 => x"69",
   785 => x"6e",
   786 => x"69",
   787 => x"74",
   788 => x"20",
   789 => x"25",
   790 => x"64",
   791 => x"0a",
   792 => x"20",
   793 => x"20",
   794 => x"00",
   795 => x"43",
   796 => x"6d",
   797 => x"64",
   798 => x"5f",
   799 => x"69",
   800 => x"6e",
   801 => x"69",
   802 => x"74",
   803 => x"0a",
   804 => x"00",
   805 => x"43",
   806 => x"4d",
   807 => x"44",
   808 => x"38",
   809 => x"5f",
   810 => x"34",
   811 => x"20",
   812 => x"72",
   813 => x"65",
   814 => x"73",
   815 => x"70",
   816 => x"6f",
   817 => x"6e",
   818 => x"73",
   819 => x"65",
   820 => x"3a",
   821 => x"20",
   822 => x"25",
   823 => x"64",
   824 => x"0a",
   825 => x"00",
   826 => x"43",
   827 => x"4d",
   828 => x"44",
   829 => x"35",
   830 => x"38",
   831 => x"20",
   832 => x"25",
   833 => x"64",
   834 => x"0a",
   835 => x"20",
   836 => x"20",
   837 => x"00",
   838 => x"43",
   839 => x"4d",
   840 => x"44",
   841 => x"35",
   842 => x"38",
   843 => x"5f",
   844 => x"32",
   845 => x"20",
   846 => x"25",
   847 => x"64",
   848 => x"0a",
   849 => x"20",
   850 => x"20",
   851 => x"00",
   852 => x"43",
   853 => x"4d",
   854 => x"44",
   855 => x"35",
   856 => x"38",
   857 => x"20",
   858 => x"25",
   859 => x"64",
   860 => x"0a",
   861 => x"20",
   862 => x"20",
   863 => x"00",
   864 => x"53",
   865 => x"44",
   866 => x"48",
   867 => x"43",
   868 => x"20",
   869 => x"49",
   870 => x"6e",
   871 => x"69",
   872 => x"74",
   873 => x"69",
   874 => x"61",
   875 => x"6c",
   876 => x"69",
   877 => x"7a",
   878 => x"61",
   879 => x"74",
   880 => x"69",
   881 => x"6f",
   882 => x"6e",
   883 => x"20",
   884 => x"65",
   885 => x"72",
   886 => x"72",
   887 => x"6f",
   888 => x"72",
   889 => x"21",
   890 => x"0a",
   891 => x"00",
   892 => x"63",
   893 => x"6d",
   894 => x"64",
   895 => x"5f",
   896 => x"43",
   897 => x"4d",
   898 => x"44",
   899 => x"38",
   900 => x"20",
   901 => x"72",
   902 => x"65",
   903 => x"73",
   904 => x"70",
   905 => x"6f",
   906 => x"6e",
   907 => x"73",
   908 => x"65",
   909 => x"3a",
   910 => x"20",
   911 => x"25",
   912 => x"64",
   913 => x"0a",
   914 => x"00",
   915 => x"52",
   916 => x"65",
   917 => x"61",
   918 => x"64",
   919 => x"20",
   920 => x"63",
   921 => x"6f",
   922 => x"6d",
   923 => x"6d",
   924 => x"61",
   925 => x"6e",
   926 => x"64",
   927 => x"20",
   928 => x"66",
   929 => x"61",
   930 => x"69",
   931 => x"6c",
   932 => x"65",
   933 => x"64",
   934 => x"20",
   935 => x"61",
   936 => x"74",
   937 => x"20",
   938 => x"25",
   939 => x"64",
   940 => x"20",
   941 => x"28",
   942 => x"25",
   943 => x"64",
   944 => x"29",
   945 => x"0a",
   946 => x"00",
   947 => x"0e",
   948 => x"5e",
   949 => x"5b",
   950 => x"5c",
   951 => x"0e",
   952 => x"c0",
   953 => x"f6",
   954 => x"e4",
   955 => x"c0",
   956 => x"c0",
   957 => x"4c",
   958 => x"c3",
   959 => x"ff",
   960 => x"97",
   961 => x"7c",
   962 => x"cc",
   963 => x"db",
   964 => x"49",
   965 => x"c0",
   966 => x"e4",
   967 => x"ee",
   968 => x"87",
   969 => x"d3",
   970 => x"4b",
   971 => x"c0",
   972 => x"1e",
   973 => x"c0",
   974 => x"ff",
   975 => x"f0",
   976 => x"c1",
   977 => x"c1",
   978 => x"49",
   979 => x"f7",
   980 => x"e1",
   981 => x"87",
   982 => x"c4",
   983 => x"86",
   984 => x"70",
   985 => x"98",
   986 => x"05",
   987 => x"c8",
   988 => x"87",
   989 => x"c3",
   990 => x"ff",
   991 => x"97",
   992 => x"7c",
   993 => x"c1",
   994 => x"48",
   995 => x"cb",
   996 => x"87",
   997 => x"fa",
   998 => x"c8",
   999 => x"87",
  1000 => x"c1",
  1001 => x"8b",
  1002 => x"05",
  1003 => x"ff",
  1004 => x"dd",
  1005 => x"87",
  1006 => x"c0",
  1007 => x"48",
  1008 => x"f9",
  1009 => x"f7",
  1010 => x"87",
  1011 => x"0e",
  1012 => x"5e",
  1013 => x"5b",
  1014 => x"5c",
  1015 => x"0e",
  1016 => x"1e",
  1017 => x"c0",
  1018 => x"f6",
  1019 => x"e4",
  1020 => x"c0",
  1021 => x"c0",
  1022 => x"4c",
  1023 => x"f9",
  1024 => x"ee",
  1025 => x"87",
  1026 => x"c6",
  1027 => x"ea",
  1028 => x"1e",
  1029 => x"c0",
  1030 => x"e1",
  1031 => x"f0",
  1032 => x"c1",
  1033 => x"c8",
  1034 => x"49",
  1035 => x"f6",
  1036 => x"e9",
  1037 => x"87",
  1038 => x"70",
  1039 => x"4b",
  1040 => x"73",
  1041 => x"1e",
  1042 => x"cd",
  1043 => x"fc",
  1044 => x"49",
  1045 => x"c0",
  1046 => x"f0",
  1047 => x"ee",
  1048 => x"87",
  1049 => x"c8",
  1050 => x"86",
  1051 => x"c1",
  1052 => x"ab",
  1053 => x"02",
  1054 => x"c8",
  1055 => x"87",
  1056 => x"fe",
  1057 => x"d0",
  1058 => x"87",
  1059 => x"c0",
  1060 => x"48",
  1061 => x"c1",
  1062 => x"f0",
  1063 => x"87",
  1064 => x"f4",
  1065 => x"e9",
  1066 => x"87",
  1067 => x"70",
  1068 => x"49",
  1069 => x"cf",
  1070 => x"ff",
  1071 => x"ff",
  1072 => x"99",
  1073 => x"c6",
  1074 => x"ea",
  1075 => x"a9",
  1076 => x"02",
  1077 => x"c8",
  1078 => x"87",
  1079 => x"fd",
  1080 => x"f9",
  1081 => x"87",
  1082 => x"c0",
  1083 => x"48",
  1084 => x"c1",
  1085 => x"d9",
  1086 => x"87",
  1087 => x"c3",
  1088 => x"ff",
  1089 => x"97",
  1090 => x"7c",
  1091 => x"c0",
  1092 => x"f1",
  1093 => x"4b",
  1094 => x"f8",
  1095 => x"fe",
  1096 => x"87",
  1097 => x"70",
  1098 => x"98",
  1099 => x"02",
  1100 => x"c0",
  1101 => x"f8",
  1102 => x"87",
  1103 => x"c0",
  1104 => x"1e",
  1105 => x"c0",
  1106 => x"ff",
  1107 => x"f0",
  1108 => x"c1",
  1109 => x"fa",
  1110 => x"49",
  1111 => x"f5",
  1112 => x"dd",
  1113 => x"87",
  1114 => x"c4",
  1115 => x"86",
  1116 => x"70",
  1117 => x"98",
  1118 => x"05",
  1119 => x"c0",
  1120 => x"e5",
  1121 => x"87",
  1122 => x"c3",
  1123 => x"ff",
  1124 => x"97",
  1125 => x"7c",
  1126 => x"97",
  1127 => x"6c",
  1128 => x"48",
  1129 => x"c4",
  1130 => x"a6",
  1131 => x"58",
  1132 => x"6e",
  1133 => x"49",
  1134 => x"c3",
  1135 => x"ff",
  1136 => x"99",
  1137 => x"97",
  1138 => x"7c",
  1139 => x"97",
  1140 => x"7c",
  1141 => x"97",
  1142 => x"7c",
  1143 => x"97",
  1144 => x"7c",
  1145 => x"c1",
  1146 => x"c0",
  1147 => x"99",
  1148 => x"02",
  1149 => x"c4",
  1150 => x"87",
  1151 => x"c1",
  1152 => x"48",
  1153 => x"d5",
  1154 => x"87",
  1155 => x"c0",
  1156 => x"48",
  1157 => x"d1",
  1158 => x"87",
  1159 => x"c2",
  1160 => x"ab",
  1161 => x"05",
  1162 => x"c4",
  1163 => x"87",
  1164 => x"c0",
  1165 => x"48",
  1166 => x"c8",
  1167 => x"87",
  1168 => x"c1",
  1169 => x"8b",
  1170 => x"05",
  1171 => x"fe",
  1172 => x"f0",
  1173 => x"87",
  1174 => x"c0",
  1175 => x"48",
  1176 => x"26",
  1177 => x"f7",
  1178 => x"ce",
  1179 => x"87",
  1180 => x"0e",
  1181 => x"5e",
  1182 => x"5b",
  1183 => x"5c",
  1184 => x"5d",
  1185 => x"0e",
  1186 => x"c0",
  1187 => x"f6",
  1188 => x"e4",
  1189 => x"c0",
  1190 => x"c0",
  1191 => x"4c",
  1192 => x"48",
  1193 => x"c4",
  1194 => x"a0",
  1195 => x"4b",
  1196 => x"c1",
  1197 => x"c3",
  1198 => x"c0",
  1199 => x"48",
  1200 => x"c1",
  1201 => x"78",
  1202 => x"c0",
  1203 => x"f6",
  1204 => x"e4",
  1205 => x"c0",
  1206 => x"c8",
  1207 => x"48",
  1208 => x"c3",
  1209 => x"ef",
  1210 => x"50",
  1211 => x"c7",
  1212 => x"4d",
  1213 => x"c3",
  1214 => x"97",
  1215 => x"7b",
  1216 => x"f6",
  1217 => x"ed",
  1218 => x"87",
  1219 => x"c2",
  1220 => x"97",
  1221 => x"7b",
  1222 => x"c3",
  1223 => x"ff",
  1224 => x"97",
  1225 => x"7c",
  1226 => x"c0",
  1227 => x"1e",
  1228 => x"c0",
  1229 => x"e5",
  1230 => x"d0",
  1231 => x"c1",
  1232 => x"c0",
  1233 => x"49",
  1234 => x"f3",
  1235 => x"e2",
  1236 => x"87",
  1237 => x"c4",
  1238 => x"86",
  1239 => x"c1",
  1240 => x"a8",
  1241 => x"05",
  1242 => x"c2",
  1243 => x"87",
  1244 => x"c1",
  1245 => x"4d",
  1246 => x"c2",
  1247 => x"ad",
  1248 => x"05",
  1249 => x"c5",
  1250 => x"87",
  1251 => x"c0",
  1252 => x"48",
  1253 => x"c0",
  1254 => x"ec",
  1255 => x"87",
  1256 => x"c1",
  1257 => x"8d",
  1258 => x"05",
  1259 => x"ff",
  1260 => x"cf",
  1261 => x"87",
  1262 => x"fc",
  1263 => x"c2",
  1264 => x"87",
  1265 => x"c1",
  1266 => x"c3",
  1267 => x"c4",
  1268 => x"58",
  1269 => x"c1",
  1270 => x"c3",
  1271 => x"c0",
  1272 => x"bf",
  1273 => x"05",
  1274 => x"cd",
  1275 => x"87",
  1276 => x"c1",
  1277 => x"1e",
  1278 => x"c0",
  1279 => x"ff",
  1280 => x"f0",
  1281 => x"c1",
  1282 => x"d0",
  1283 => x"49",
  1284 => x"f2",
  1285 => x"f0",
  1286 => x"87",
  1287 => x"c4",
  1288 => x"86",
  1289 => x"c3",
  1290 => x"ff",
  1291 => x"97",
  1292 => x"7c",
  1293 => x"c3",
  1294 => x"53",
  1295 => x"c3",
  1296 => x"ff",
  1297 => x"54",
  1298 => x"c1",
  1299 => x"48",
  1300 => x"f5",
  1301 => x"d1",
  1302 => x"87",
  1303 => x"0e",
  1304 => x"5e",
  1305 => x"5b",
  1306 => x"5c",
  1307 => x"5d",
  1308 => x"0e",
  1309 => x"f8",
  1310 => x"86",
  1311 => x"71",
  1312 => x"4a",
  1313 => x"c0",
  1314 => x"f6",
  1315 => x"e4",
  1316 => x"c0",
  1317 => x"c0",
  1318 => x"4b",
  1319 => x"c0",
  1320 => x"7e",
  1321 => x"c3",
  1322 => x"ff",
  1323 => x"97",
  1324 => x"7b",
  1325 => x"c0",
  1326 => x"f6",
  1327 => x"e4",
  1328 => x"c0",
  1329 => x"c4",
  1330 => x"48",
  1331 => x"c2",
  1332 => x"50",
  1333 => x"c0",
  1334 => x"f6",
  1335 => x"e4",
  1336 => x"c0",
  1337 => x"c8",
  1338 => x"48",
  1339 => x"c7",
  1340 => x"50",
  1341 => x"c3",
  1342 => x"ff",
  1343 => x"97",
  1344 => x"7b",
  1345 => x"72",
  1346 => x"1e",
  1347 => x"c0",
  1348 => x"ff",
  1349 => x"f0",
  1350 => x"c1",
  1351 => x"d1",
  1352 => x"49",
  1353 => x"f1",
  1354 => x"eb",
  1355 => x"87",
  1356 => x"c4",
  1357 => x"86",
  1358 => x"70",
  1359 => x"98",
  1360 => x"05",
  1361 => x"c1",
  1362 => x"ca",
  1363 => x"87",
  1364 => x"c5",
  1365 => x"ee",
  1366 => x"cd",
  1367 => x"df",
  1368 => x"4c",
  1369 => x"c3",
  1370 => x"ff",
  1371 => x"97",
  1372 => x"7b",
  1373 => x"97",
  1374 => x"6b",
  1375 => x"48",
  1376 => x"c8",
  1377 => x"a6",
  1378 => x"58",
  1379 => x"c4",
  1380 => x"66",
  1381 => x"49",
  1382 => x"c3",
  1383 => x"ff",
  1384 => x"99",
  1385 => x"c3",
  1386 => x"fe",
  1387 => x"a9",
  1388 => x"05",
  1389 => x"de",
  1390 => x"87",
  1391 => x"c0",
  1392 => x"4d",
  1393 => x"ef",
  1394 => x"e0",
  1395 => x"87",
  1396 => x"d8",
  1397 => x"66",
  1398 => x"08",
  1399 => x"78",
  1400 => x"08",
  1401 => x"d8",
  1402 => x"66",
  1403 => x"48",
  1404 => x"c4",
  1405 => x"80",
  1406 => x"dc",
  1407 => x"a6",
  1408 => x"58",
  1409 => x"c1",
  1410 => x"85",
  1411 => x"c2",
  1412 => x"c0",
  1413 => x"b7",
  1414 => x"ad",
  1415 => x"04",
  1416 => x"e7",
  1417 => x"87",
  1418 => x"c1",
  1419 => x"4c",
  1420 => x"7e",
  1421 => x"c1",
  1422 => x"8c",
  1423 => x"05",
  1424 => x"ff",
  1425 => x"c6",
  1426 => x"87",
  1427 => x"c3",
  1428 => x"ff",
  1429 => x"53",
  1430 => x"c0",
  1431 => x"f6",
  1432 => x"e4",
  1433 => x"c0",
  1434 => x"c4",
  1435 => x"48",
  1436 => x"c3",
  1437 => x"50",
  1438 => x"6e",
  1439 => x"48",
  1440 => x"f8",
  1441 => x"8e",
  1442 => x"f3",
  1443 => x"c3",
  1444 => x"87",
  1445 => x"1e",
  1446 => x"73",
  1447 => x"1e",
  1448 => x"71",
  1449 => x"4b",
  1450 => x"73",
  1451 => x"49",
  1452 => x"d8",
  1453 => x"29",
  1454 => x"c3",
  1455 => x"ff",
  1456 => x"99",
  1457 => x"73",
  1458 => x"4a",
  1459 => x"c8",
  1460 => x"2a",
  1461 => x"cf",
  1462 => x"fc",
  1463 => x"c0",
  1464 => x"9a",
  1465 => x"72",
  1466 => x"b1",
  1467 => x"73",
  1468 => x"4a",
  1469 => x"c8",
  1470 => x"32",
  1471 => x"c0",
  1472 => x"ff",
  1473 => x"f0",
  1474 => x"c0",
  1475 => x"c0",
  1476 => x"9a",
  1477 => x"72",
  1478 => x"b1",
  1479 => x"73",
  1480 => x"4a",
  1481 => x"d8",
  1482 => x"32",
  1483 => x"ff",
  1484 => x"c0",
  1485 => x"c0",
  1486 => x"c0",
  1487 => x"c0",
  1488 => x"9a",
  1489 => x"72",
  1490 => x"b1",
  1491 => x"71",
  1492 => x"48",
  1493 => x"c4",
  1494 => x"87",
  1495 => x"26",
  1496 => x"4d",
  1497 => x"26",
  1498 => x"4c",
  1499 => x"26",
  1500 => x"4b",
  1501 => x"26",
  1502 => x"4f",
  1503 => x"1e",
  1504 => x"73",
  1505 => x"1e",
  1506 => x"71",
  1507 => x"4b",
  1508 => x"73",
  1509 => x"49",
  1510 => x"c8",
  1511 => x"29",
  1512 => x"c3",
  1513 => x"ff",
  1514 => x"99",
  1515 => x"73",
  1516 => x"4a",
  1517 => x"c8",
  1518 => x"32",
  1519 => x"cf",
  1520 => x"fc",
  1521 => x"c0",
  1522 => x"9a",
  1523 => x"72",
  1524 => x"b1",
  1525 => x"71",
  1526 => x"48",
  1527 => x"e2",
  1528 => x"87",
  1529 => x"0e",
  1530 => x"5e",
  1531 => x"5b",
  1532 => x"5c",
  1533 => x"0e",
  1534 => x"71",
  1535 => x"4b",
  1536 => x"c0",
  1537 => x"4c",
  1538 => x"d0",
  1539 => x"66",
  1540 => x"48",
  1541 => x"c0",
  1542 => x"b7",
  1543 => x"a8",
  1544 => x"06",
  1545 => x"c0",
  1546 => x"e3",
  1547 => x"87",
  1548 => x"13",
  1549 => x"4a",
  1550 => x"cc",
  1551 => x"66",
  1552 => x"97",
  1553 => x"bf",
  1554 => x"49",
  1555 => x"cc",
  1556 => x"66",
  1557 => x"48",
  1558 => x"c1",
  1559 => x"80",
  1560 => x"d0",
  1561 => x"a6",
  1562 => x"58",
  1563 => x"71",
  1564 => x"b7",
  1565 => x"aa",
  1566 => x"02",
  1567 => x"c4",
  1568 => x"87",
  1569 => x"c1",
  1570 => x"48",
  1571 => x"cc",
  1572 => x"87",
  1573 => x"c1",
  1574 => x"84",
  1575 => x"d0",
  1576 => x"66",
  1577 => x"b7",
  1578 => x"ac",
  1579 => x"04",
  1580 => x"ff",
  1581 => x"dd",
  1582 => x"87",
  1583 => x"c0",
  1584 => x"48",
  1585 => x"c2",
  1586 => x"87",
  1587 => x"26",
  1588 => x"4d",
  1589 => x"26",
  1590 => x"4c",
  1591 => x"26",
  1592 => x"4b",
  1593 => x"26",
  1594 => x"4f",
  1595 => x"0e",
  1596 => x"5e",
  1597 => x"5b",
  1598 => x"5c",
  1599 => x"5d",
  1600 => x"0e",
  1601 => x"c1",
  1602 => x"cc",
  1603 => x"c2",
  1604 => x"48",
  1605 => x"ff",
  1606 => x"78",
  1607 => x"c1",
  1608 => x"cb",
  1609 => x"d2",
  1610 => x"48",
  1611 => x"c0",
  1612 => x"78",
  1613 => x"c0",
  1614 => x"e6",
  1615 => x"f0",
  1616 => x"49",
  1617 => x"da",
  1618 => x"e3",
  1619 => x"87",
  1620 => x"c1",
  1621 => x"c3",
  1622 => x"ca",
  1623 => x"1e",
  1624 => x"c0",
  1625 => x"49",
  1626 => x"fa",
  1627 => x"fa",
  1628 => x"87",
  1629 => x"c4",
  1630 => x"86",
  1631 => x"70",
  1632 => x"98",
  1633 => x"05",
  1634 => x"c5",
  1635 => x"87",
  1636 => x"c0",
  1637 => x"48",
  1638 => x"cb",
  1639 => x"c1",
  1640 => x"87",
  1641 => x"c0",
  1642 => x"4b",
  1643 => x"c1",
  1644 => x"cb",
  1645 => x"fe",
  1646 => x"48",
  1647 => x"c1",
  1648 => x"78",
  1649 => x"c8",
  1650 => x"1e",
  1651 => x"c0",
  1652 => x"e6",
  1653 => x"fd",
  1654 => x"1e",
  1655 => x"c1",
  1656 => x"c4",
  1657 => x"c0",
  1658 => x"49",
  1659 => x"fd",
  1660 => x"fb",
  1661 => x"87",
  1662 => x"c8",
  1663 => x"86",
  1664 => x"70",
  1665 => x"98",
  1666 => x"05",
  1667 => x"c6",
  1668 => x"87",
  1669 => x"c1",
  1670 => x"cb",
  1671 => x"fe",
  1672 => x"48",
  1673 => x"c0",
  1674 => x"78",
  1675 => x"c8",
  1676 => x"1e",
  1677 => x"c0",
  1678 => x"e7",
  1679 => x"c6",
  1680 => x"1e",
  1681 => x"c1",
  1682 => x"c4",
  1683 => x"dc",
  1684 => x"49",
  1685 => x"fd",
  1686 => x"e1",
  1687 => x"87",
  1688 => x"c8",
  1689 => x"86",
  1690 => x"70",
  1691 => x"98",
  1692 => x"05",
  1693 => x"c6",
  1694 => x"87",
  1695 => x"c1",
  1696 => x"cb",
  1697 => x"fe",
  1698 => x"48",
  1699 => x"c0",
  1700 => x"78",
  1701 => x"c8",
  1702 => x"1e",
  1703 => x"c0",
  1704 => x"e7",
  1705 => x"cf",
  1706 => x"1e",
  1707 => x"c1",
  1708 => x"c4",
  1709 => x"dc",
  1710 => x"49",
  1711 => x"fd",
  1712 => x"c7",
  1713 => x"87",
  1714 => x"c8",
  1715 => x"86",
  1716 => x"70",
  1717 => x"98",
  1718 => x"05",
  1719 => x"c5",
  1720 => x"87",
  1721 => x"c0",
  1722 => x"48",
  1723 => x"c9",
  1724 => x"ec",
  1725 => x"87",
  1726 => x"c1",
  1727 => x"cb",
  1728 => x"fe",
  1729 => x"bf",
  1730 => x"1e",
  1731 => x"c0",
  1732 => x"e7",
  1733 => x"d8",
  1734 => x"1e",
  1735 => x"c0",
  1736 => x"e5",
  1737 => x"fc",
  1738 => x"87",
  1739 => x"c8",
  1740 => x"86",
  1741 => x"c1",
  1742 => x"cb",
  1743 => x"fe",
  1744 => x"bf",
  1745 => x"02",
  1746 => x"c1",
  1747 => x"f4",
  1748 => x"87",
  1749 => x"c1",
  1750 => x"c3",
  1751 => x"ca",
  1752 => x"4d",
  1753 => x"48",
  1754 => x"c6",
  1755 => x"fe",
  1756 => x"a0",
  1757 => x"4c",
  1758 => x"c8",
  1759 => x"c0",
  1760 => x"1e",
  1761 => x"70",
  1762 => x"49",
  1763 => x"d8",
  1764 => x"fb",
  1765 => x"87",
  1766 => x"c4",
  1767 => x"86",
  1768 => x"c8",
  1769 => x"a4",
  1770 => x"49",
  1771 => x"69",
  1772 => x"4b",
  1773 => x"c1",
  1774 => x"cb",
  1775 => x"c8",
  1776 => x"9f",
  1777 => x"bf",
  1778 => x"49",
  1779 => x"c5",
  1780 => x"d6",
  1781 => x"ea",
  1782 => x"a9",
  1783 => x"05",
  1784 => x"c0",
  1785 => x"cc",
  1786 => x"87",
  1787 => x"c8",
  1788 => x"a4",
  1789 => x"4a",
  1790 => x"6a",
  1791 => x"49",
  1792 => x"fa",
  1793 => x"e2",
  1794 => x"87",
  1795 => x"70",
  1796 => x"4b",
  1797 => x"db",
  1798 => x"87",
  1799 => x"c7",
  1800 => x"fe",
  1801 => x"a5",
  1802 => x"49",
  1803 => x"9f",
  1804 => x"69",
  1805 => x"49",
  1806 => x"ca",
  1807 => x"e9",
  1808 => x"d5",
  1809 => x"a9",
  1810 => x"02",
  1811 => x"c0",
  1812 => x"cc",
  1813 => x"87",
  1814 => x"c0",
  1815 => x"e4",
  1816 => x"ed",
  1817 => x"49",
  1818 => x"d7",
  1819 => x"da",
  1820 => x"87",
  1821 => x"c0",
  1822 => x"48",
  1823 => x"c8",
  1824 => x"c8",
  1825 => x"87",
  1826 => x"73",
  1827 => x"1e",
  1828 => x"c0",
  1829 => x"e5",
  1830 => x"cb",
  1831 => x"1e",
  1832 => x"c0",
  1833 => x"e4",
  1834 => x"db",
  1835 => x"87",
  1836 => x"c1",
  1837 => x"c3",
  1838 => x"ca",
  1839 => x"1e",
  1840 => x"73",
  1841 => x"49",
  1842 => x"f7",
  1843 => x"e2",
  1844 => x"87",
  1845 => x"cc",
  1846 => x"86",
  1847 => x"70",
  1848 => x"98",
  1849 => x"05",
  1850 => x"c0",
  1851 => x"c5",
  1852 => x"87",
  1853 => x"c0",
  1854 => x"48",
  1855 => x"c7",
  1856 => x"e8",
  1857 => x"87",
  1858 => x"c0",
  1859 => x"e5",
  1860 => x"e3",
  1861 => x"49",
  1862 => x"d6",
  1863 => x"ee",
  1864 => x"87",
  1865 => x"c8",
  1866 => x"c0",
  1867 => x"1e",
  1868 => x"c1",
  1869 => x"c3",
  1870 => x"ca",
  1871 => x"49",
  1872 => x"d7",
  1873 => x"ce",
  1874 => x"87",
  1875 => x"c0",
  1876 => x"e7",
  1877 => x"eb",
  1878 => x"1e",
  1879 => x"c0",
  1880 => x"e3",
  1881 => x"ec",
  1882 => x"87",
  1883 => x"c8",
  1884 => x"1e",
  1885 => x"c0",
  1886 => x"e8",
  1887 => x"c3",
  1888 => x"1e",
  1889 => x"c1",
  1890 => x"c4",
  1891 => x"dc",
  1892 => x"49",
  1893 => x"fa",
  1894 => x"d1",
  1895 => x"87",
  1896 => x"d0",
  1897 => x"86",
  1898 => x"70",
  1899 => x"98",
  1900 => x"05",
  1901 => x"c0",
  1902 => x"c9",
  1903 => x"87",
  1904 => x"c1",
  1905 => x"cb",
  1906 => x"d2",
  1907 => x"48",
  1908 => x"c1",
  1909 => x"78",
  1910 => x"c0",
  1911 => x"e4",
  1912 => x"87",
  1913 => x"c8",
  1914 => x"1e",
  1915 => x"c0",
  1916 => x"e8",
  1917 => x"cc",
  1918 => x"1e",
  1919 => x"c1",
  1920 => x"c4",
  1921 => x"c0",
  1922 => x"49",
  1923 => x"f9",
  1924 => x"f3",
  1925 => x"87",
  1926 => x"c8",
  1927 => x"86",
  1928 => x"70",
  1929 => x"98",
  1930 => x"02",
  1931 => x"c0",
  1932 => x"cf",
  1933 => x"87",
  1934 => x"c0",
  1935 => x"e6",
  1936 => x"ca",
  1937 => x"1e",
  1938 => x"c0",
  1939 => x"e2",
  1940 => x"f1",
  1941 => x"87",
  1942 => x"c4",
  1943 => x"86",
  1944 => x"c0",
  1945 => x"48",
  1946 => x"c6",
  1947 => x"cd",
  1948 => x"87",
  1949 => x"c1",
  1950 => x"cb",
  1951 => x"c8",
  1952 => x"97",
  1953 => x"bf",
  1954 => x"49",
  1955 => x"c1",
  1956 => x"d5",
  1957 => x"a9",
  1958 => x"05",
  1959 => x"c0",
  1960 => x"cd",
  1961 => x"87",
  1962 => x"c1",
  1963 => x"cb",
  1964 => x"c9",
  1965 => x"97",
  1966 => x"bf",
  1967 => x"49",
  1968 => x"c2",
  1969 => x"ea",
  1970 => x"a9",
  1971 => x"02",
  1972 => x"c0",
  1973 => x"c5",
  1974 => x"87",
  1975 => x"c0",
  1976 => x"48",
  1977 => x"c5",
  1978 => x"ee",
  1979 => x"87",
  1980 => x"c1",
  1981 => x"c3",
  1982 => x"ca",
  1983 => x"97",
  1984 => x"bf",
  1985 => x"49",
  1986 => x"c3",
  1987 => x"e9",
  1988 => x"a9",
  1989 => x"02",
  1990 => x"c0",
  1991 => x"d2",
  1992 => x"87",
  1993 => x"c1",
  1994 => x"c3",
  1995 => x"ca",
  1996 => x"97",
  1997 => x"bf",
  1998 => x"49",
  1999 => x"c3",
  2000 => x"eb",
  2001 => x"a9",
  2002 => x"02",
  2003 => x"c0",
  2004 => x"c5",
  2005 => x"87",
  2006 => x"c0",
  2007 => x"48",
  2008 => x"c5",
  2009 => x"cf",
  2010 => x"87",
  2011 => x"c1",
  2012 => x"c3",
  2013 => x"d5",
  2014 => x"97",
  2015 => x"bf",
  2016 => x"49",
  2017 => x"71",
  2018 => x"99",
  2019 => x"05",
  2020 => x"c0",
  2021 => x"cc",
  2022 => x"87",
  2023 => x"c1",
  2024 => x"c3",
  2025 => x"d6",
  2026 => x"97",
  2027 => x"bf",
  2028 => x"49",
  2029 => x"c2",
  2030 => x"a9",
  2031 => x"02",
  2032 => x"c0",
  2033 => x"c5",
  2034 => x"87",
  2035 => x"c0",
  2036 => x"48",
  2037 => x"c4",
  2038 => x"f2",
  2039 => x"87",
  2040 => x"c1",
  2041 => x"c3",
  2042 => x"d7",
  2043 => x"97",
  2044 => x"bf",
  2045 => x"48",
  2046 => x"c1",
  2047 => x"cb",
  2048 => x"ce",
  2049 => x"58",
  2050 => x"c1",
  2051 => x"cb",
  2052 => x"ca",
  2053 => x"bf",
  2054 => x"48",
  2055 => x"c1",
  2056 => x"88",
  2057 => x"c1",
  2058 => x"cb",
  2059 => x"d2",
  2060 => x"58",
  2061 => x"c1",
  2062 => x"c3",
  2063 => x"d8",
  2064 => x"97",
  2065 => x"bf",
  2066 => x"49",
  2067 => x"73",
  2068 => x"81",
  2069 => x"c1",
  2070 => x"c3",
  2071 => x"d9",
  2072 => x"97",
  2073 => x"bf",
  2074 => x"4a",
  2075 => x"c8",
  2076 => x"32",
  2077 => x"c1",
  2078 => x"cb",
  2079 => x"de",
  2080 => x"48",
  2081 => x"72",
  2082 => x"a1",
  2083 => x"78",
  2084 => x"c1",
  2085 => x"c3",
  2086 => x"da",
  2087 => x"97",
  2088 => x"bf",
  2089 => x"48",
  2090 => x"c1",
  2091 => x"cb",
  2092 => x"f6",
  2093 => x"58",
  2094 => x"c1",
  2095 => x"cb",
  2096 => x"d2",
  2097 => x"bf",
  2098 => x"02",
  2099 => x"c2",
  2100 => x"e2",
  2101 => x"87",
  2102 => x"c8",
  2103 => x"1e",
  2104 => x"c0",
  2105 => x"e6",
  2106 => x"e7",
  2107 => x"1e",
  2108 => x"c1",
  2109 => x"c4",
  2110 => x"dc",
  2111 => x"49",
  2112 => x"f6",
  2113 => x"f6",
  2114 => x"87",
  2115 => x"c8",
  2116 => x"86",
  2117 => x"70",
  2118 => x"98",
  2119 => x"02",
  2120 => x"c0",
  2121 => x"c5",
  2122 => x"87",
  2123 => x"c0",
  2124 => x"48",
  2125 => x"c3",
  2126 => x"da",
  2127 => x"87",
  2128 => x"c1",
  2129 => x"cb",
  2130 => x"ca",
  2131 => x"bf",
  2132 => x"48",
  2133 => x"c4",
  2134 => x"30",
  2135 => x"c1",
  2136 => x"cb",
  2137 => x"fa",
  2138 => x"58",
  2139 => x"c1",
  2140 => x"cb",
  2141 => x"ca",
  2142 => x"bf",
  2143 => x"4a",
  2144 => x"c1",
  2145 => x"cb",
  2146 => x"f2",
  2147 => x"5a",
  2148 => x"c1",
  2149 => x"c3",
  2150 => x"ef",
  2151 => x"97",
  2152 => x"bf",
  2153 => x"49",
  2154 => x"c8",
  2155 => x"31",
  2156 => x"c1",
  2157 => x"c3",
  2158 => x"ee",
  2159 => x"97",
  2160 => x"bf",
  2161 => x"4b",
  2162 => x"73",
  2163 => x"a1",
  2164 => x"49",
  2165 => x"c1",
  2166 => x"c3",
  2167 => x"f0",
  2168 => x"97",
  2169 => x"bf",
  2170 => x"4b",
  2171 => x"d0",
  2172 => x"33",
  2173 => x"73",
  2174 => x"a1",
  2175 => x"49",
  2176 => x"c1",
  2177 => x"c3",
  2178 => x"f1",
  2179 => x"97",
  2180 => x"bf",
  2181 => x"4b",
  2182 => x"d8",
  2183 => x"33",
  2184 => x"73",
  2185 => x"a1",
  2186 => x"49",
  2187 => x"c1",
  2188 => x"cb",
  2189 => x"fe",
  2190 => x"59",
  2191 => x"c1",
  2192 => x"cb",
  2193 => x"f2",
  2194 => x"bf",
  2195 => x"91",
  2196 => x"c1",
  2197 => x"cb",
  2198 => x"de",
  2199 => x"bf",
  2200 => x"81",
  2201 => x"c1",
  2202 => x"cb",
  2203 => x"e6",
  2204 => x"59",
  2205 => x"c1",
  2206 => x"c3",
  2207 => x"f7",
  2208 => x"97",
  2209 => x"bf",
  2210 => x"4b",
  2211 => x"c8",
  2212 => x"33",
  2213 => x"c1",
  2214 => x"c3",
  2215 => x"f6",
  2216 => x"97",
  2217 => x"bf",
  2218 => x"4c",
  2219 => x"74",
  2220 => x"a3",
  2221 => x"4b",
  2222 => x"c1",
  2223 => x"c3",
  2224 => x"f8",
  2225 => x"97",
  2226 => x"bf",
  2227 => x"4c",
  2228 => x"d0",
  2229 => x"34",
  2230 => x"74",
  2231 => x"a3",
  2232 => x"4b",
  2233 => x"c1",
  2234 => x"c3",
  2235 => x"f9",
  2236 => x"97",
  2237 => x"bf",
  2238 => x"4c",
  2239 => x"cf",
  2240 => x"9c",
  2241 => x"d8",
  2242 => x"34",
  2243 => x"74",
  2244 => x"a3",
  2245 => x"4b",
  2246 => x"c1",
  2247 => x"cb",
  2248 => x"ea",
  2249 => x"5b",
  2250 => x"c2",
  2251 => x"8b",
  2252 => x"73",
  2253 => x"92",
  2254 => x"c1",
  2255 => x"cb",
  2256 => x"ea",
  2257 => x"48",
  2258 => x"72",
  2259 => x"a1",
  2260 => x"78",
  2261 => x"c1",
  2262 => x"d0",
  2263 => x"87",
  2264 => x"c1",
  2265 => x"c3",
  2266 => x"dc",
  2267 => x"97",
  2268 => x"bf",
  2269 => x"49",
  2270 => x"c8",
  2271 => x"31",
  2272 => x"c1",
  2273 => x"c3",
  2274 => x"db",
  2275 => x"97",
  2276 => x"bf",
  2277 => x"4a",
  2278 => x"72",
  2279 => x"a1",
  2280 => x"49",
  2281 => x"c1",
  2282 => x"cb",
  2283 => x"fa",
  2284 => x"59",
  2285 => x"c5",
  2286 => x"31",
  2287 => x"c7",
  2288 => x"ff",
  2289 => x"81",
  2290 => x"c9",
  2291 => x"29",
  2292 => x"c1",
  2293 => x"cb",
  2294 => x"f2",
  2295 => x"59",
  2296 => x"c1",
  2297 => x"c3",
  2298 => x"e1",
  2299 => x"97",
  2300 => x"bf",
  2301 => x"4a",
  2302 => x"c8",
  2303 => x"32",
  2304 => x"c1",
  2305 => x"c3",
  2306 => x"e0",
  2307 => x"97",
  2308 => x"bf",
  2309 => x"4b",
  2310 => x"73",
  2311 => x"a2",
  2312 => x"4a",
  2313 => x"c1",
  2314 => x"cb",
  2315 => x"fe",
  2316 => x"5a",
  2317 => x"c1",
  2318 => x"cb",
  2319 => x"f2",
  2320 => x"bf",
  2321 => x"92",
  2322 => x"c1",
  2323 => x"cb",
  2324 => x"de",
  2325 => x"bf",
  2326 => x"82",
  2327 => x"c1",
  2328 => x"cb",
  2329 => x"ee",
  2330 => x"5a",
  2331 => x"c1",
  2332 => x"cb",
  2333 => x"e6",
  2334 => x"48",
  2335 => x"c0",
  2336 => x"78",
  2337 => x"c1",
  2338 => x"cb",
  2339 => x"e2",
  2340 => x"48",
  2341 => x"72",
  2342 => x"a1",
  2343 => x"78",
  2344 => x"c1",
  2345 => x"48",
  2346 => x"f4",
  2347 => x"c6",
  2348 => x"87",
  2349 => x"4e",
  2350 => x"6f",
  2351 => x"20",
  2352 => x"70",
  2353 => x"61",
  2354 => x"72",
  2355 => x"74",
  2356 => x"69",
  2357 => x"74",
  2358 => x"69",
  2359 => x"6f",
  2360 => x"6e",
  2361 => x"20",
  2362 => x"73",
  2363 => x"69",
  2364 => x"67",
  2365 => x"6e",
  2366 => x"61",
  2367 => x"74",
  2368 => x"75",
  2369 => x"72",
  2370 => x"65",
  2371 => x"20",
  2372 => x"66",
  2373 => x"6f",
  2374 => x"75",
  2375 => x"6e",
  2376 => x"64",
  2377 => x"0a",
  2378 => x"00",
  2379 => x"52",
  2380 => x"65",
  2381 => x"61",
  2382 => x"64",
  2383 => x"69",
  2384 => x"6e",
  2385 => x"67",
  2386 => x"20",
  2387 => x"62",
  2388 => x"6f",
  2389 => x"6f",
  2390 => x"74",
  2391 => x"20",
  2392 => x"73",
  2393 => x"65",
  2394 => x"63",
  2395 => x"74",
  2396 => x"6f",
  2397 => x"72",
  2398 => x"20",
  2399 => x"25",
  2400 => x"64",
  2401 => x"0a",
  2402 => x"00",
  2403 => x"52",
  2404 => x"65",
  2405 => x"61",
  2406 => x"64",
  2407 => x"20",
  2408 => x"62",
  2409 => x"6f",
  2410 => x"6f",
  2411 => x"74",
  2412 => x"20",
  2413 => x"73",
  2414 => x"65",
  2415 => x"63",
  2416 => x"74",
  2417 => x"6f",
  2418 => x"72",
  2419 => x"20",
  2420 => x"66",
  2421 => x"72",
  2422 => x"6f",
  2423 => x"6d",
  2424 => x"20",
  2425 => x"66",
  2426 => x"69",
  2427 => x"72",
  2428 => x"73",
  2429 => x"74",
  2430 => x"20",
  2431 => x"70",
  2432 => x"61",
  2433 => x"72",
  2434 => x"74",
  2435 => x"69",
  2436 => x"74",
  2437 => x"69",
  2438 => x"6f",
  2439 => x"6e",
  2440 => x"0a",
  2441 => x"00",
  2442 => x"55",
  2443 => x"6e",
  2444 => x"73",
  2445 => x"75",
  2446 => x"70",
  2447 => x"70",
  2448 => x"6f",
  2449 => x"72",
  2450 => x"74",
  2451 => x"65",
  2452 => x"64",
  2453 => x"20",
  2454 => x"70",
  2455 => x"61",
  2456 => x"72",
  2457 => x"74",
  2458 => x"69",
  2459 => x"74",
  2460 => x"69",
  2461 => x"6f",
  2462 => x"6e",
  2463 => x"20",
  2464 => x"74",
  2465 => x"79",
  2466 => x"70",
  2467 => x"65",
  2468 => x"21",
  2469 => x"0d",
  2470 => x"00",
  2471 => x"46",
  2472 => x"41",
  2473 => x"54",
  2474 => x"33",
  2475 => x"32",
  2476 => x"20",
  2477 => x"20",
  2478 => x"20",
  2479 => x"00",
  2480 => x"52",
  2481 => x"65",
  2482 => x"61",
  2483 => x"64",
  2484 => x"69",
  2485 => x"6e",
  2486 => x"67",
  2487 => x"20",
  2488 => x"4d",
  2489 => x"42",
  2490 => x"52",
  2491 => x"0a",
  2492 => x"00",
  2493 => x"46",
  2494 => x"41",
  2495 => x"54",
  2496 => x"31",
  2497 => x"36",
  2498 => x"20",
  2499 => x"20",
  2500 => x"20",
  2501 => x"00",
  2502 => x"46",
  2503 => x"41",
  2504 => x"54",
  2505 => x"33",
  2506 => x"32",
  2507 => x"20",
  2508 => x"20",
  2509 => x"20",
  2510 => x"00",
  2511 => x"46",
  2512 => x"41",
  2513 => x"54",
  2514 => x"31",
  2515 => x"32",
  2516 => x"20",
  2517 => x"20",
  2518 => x"20",
  2519 => x"00",
  2520 => x"50",
  2521 => x"61",
  2522 => x"72",
  2523 => x"74",
  2524 => x"69",
  2525 => x"74",
  2526 => x"69",
  2527 => x"6f",
  2528 => x"6e",
  2529 => x"63",
  2530 => x"6f",
  2531 => x"75",
  2532 => x"6e",
  2533 => x"74",
  2534 => x"20",
  2535 => x"25",
  2536 => x"64",
  2537 => x"0a",
  2538 => x"00",
  2539 => x"48",
  2540 => x"75",
  2541 => x"6e",
  2542 => x"74",
  2543 => x"69",
  2544 => x"6e",
  2545 => x"67",
  2546 => x"20",
  2547 => x"66",
  2548 => x"6f",
  2549 => x"72",
  2550 => x"20",
  2551 => x"66",
  2552 => x"69",
  2553 => x"6c",
  2554 => x"65",
  2555 => x"73",
  2556 => x"79",
  2557 => x"73",
  2558 => x"74",
  2559 => x"65",
  2560 => x"6d",
  2561 => x"0a",
  2562 => x"00",
  2563 => x"46",
  2564 => x"41",
  2565 => x"54",
  2566 => x"33",
  2567 => x"32",
  2568 => x"20",
  2569 => x"20",
  2570 => x"20",
  2571 => x"00",
  2572 => x"46",
  2573 => x"41",
  2574 => x"54",
  2575 => x"31",
  2576 => x"36",
  2577 => x"20",
  2578 => x"20",
  2579 => x"20",
  2580 => x"00",
  2581 => x"52",
  2582 => x"65",
  2583 => x"61",
  2584 => x"64",
  2585 => x"69",
  2586 => x"6e",
  2587 => x"67",
  2588 => x"20",
  2589 => x"64",
  2590 => x"69",
  2591 => x"72",
  2592 => x"65",
  2593 => x"63",
  2594 => x"74",
  2595 => x"6f",
  2596 => x"72",
  2597 => x"79",
  2598 => x"20",
  2599 => x"73",
  2600 => x"65",
  2601 => x"63",
  2602 => x"74",
  2603 => x"6f",
  2604 => x"72",
  2605 => x"20",
  2606 => x"25",
  2607 => x"64",
  2608 => x"0a",
  2609 => x"00",
  2610 => x"66",
  2611 => x"69",
  2612 => x"6c",
  2613 => x"65",
  2614 => x"20",
  2615 => x"22",
  2616 => x"25",
  2617 => x"73",
  2618 => x"22",
  2619 => x"20",
  2620 => x"66",
  2621 => x"6f",
  2622 => x"75",
  2623 => x"6e",
  2624 => x"64",
  2625 => x"0d",
  2626 => x"00",
  2627 => x"47",
  2628 => x"65",
  2629 => x"74",
  2630 => x"46",
  2631 => x"41",
  2632 => x"54",
  2633 => x"4c",
  2634 => x"69",
  2635 => x"6e",
  2636 => x"6b",
  2637 => x"20",
  2638 => x"72",
  2639 => x"65",
  2640 => x"74",
  2641 => x"75",
  2642 => x"72",
  2643 => x"6e",
  2644 => x"65",
  2645 => x"64",
  2646 => x"20",
  2647 => x"25",
  2648 => x"64",
  2649 => x"0a",
  2650 => x"00",
  2651 => x"43",
  2652 => x"61",
  2653 => x"6e",
  2654 => x"27",
  2655 => x"74",
  2656 => x"20",
  2657 => x"6f",
  2658 => x"70",
  2659 => x"65",
  2660 => x"6e",
  2661 => x"20",
  2662 => x"25",
  2663 => x"73",
  2664 => x"0a",
  2665 => x"00",
  2666 => x"0e",
  2667 => x"5e",
  2668 => x"5b",
  2669 => x"5c",
  2670 => x"5d",
  2671 => x"0e",
  2672 => x"71",
  2673 => x"4a",
  2674 => x"c1",
  2675 => x"cb",
  2676 => x"d2",
  2677 => x"bf",
  2678 => x"02",
  2679 => x"cc",
  2680 => x"87",
  2681 => x"72",
  2682 => x"4b",
  2683 => x"c7",
  2684 => x"b7",
  2685 => x"2b",
  2686 => x"72",
  2687 => x"4c",
  2688 => x"c1",
  2689 => x"ff",
  2690 => x"9c",
  2691 => x"ca",
  2692 => x"87",
  2693 => x"72",
  2694 => x"4b",
  2695 => x"c8",
  2696 => x"b7",
  2697 => x"2b",
  2698 => x"72",
  2699 => x"4c",
  2700 => x"c3",
  2701 => x"ff",
  2702 => x"9c",
  2703 => x"c1",
  2704 => x"cc",
  2705 => x"c2",
  2706 => x"bf",
  2707 => x"ab",
  2708 => x"02",
  2709 => x"de",
  2710 => x"87",
  2711 => x"c1",
  2712 => x"c3",
  2713 => x"ca",
  2714 => x"1e",
  2715 => x"c1",
  2716 => x"cb",
  2717 => x"de",
  2718 => x"bf",
  2719 => x"49",
  2720 => x"73",
  2721 => x"81",
  2722 => x"e9",
  2723 => x"f2",
  2724 => x"87",
  2725 => x"c4",
  2726 => x"86",
  2727 => x"70",
  2728 => x"98",
  2729 => x"05",
  2730 => x"c5",
  2731 => x"87",
  2732 => x"c0",
  2733 => x"48",
  2734 => x"c0",
  2735 => x"f6",
  2736 => x"87",
  2737 => x"c1",
  2738 => x"cc",
  2739 => x"c6",
  2740 => x"5b",
  2741 => x"c1",
  2742 => x"cb",
  2743 => x"d2",
  2744 => x"bf",
  2745 => x"02",
  2746 => x"d9",
  2747 => x"87",
  2748 => x"74",
  2749 => x"4a",
  2750 => x"c4",
  2751 => x"92",
  2752 => x"c1",
  2753 => x"c3",
  2754 => x"ca",
  2755 => x"82",
  2756 => x"6a",
  2757 => x"49",
  2758 => x"eb",
  2759 => x"dc",
  2760 => x"87",
  2761 => x"70",
  2762 => x"49",
  2763 => x"71",
  2764 => x"4d",
  2765 => x"cf",
  2766 => x"ff",
  2767 => x"ff",
  2768 => x"ff",
  2769 => x"ff",
  2770 => x"9d",
  2771 => x"d0",
  2772 => x"87",
  2773 => x"74",
  2774 => x"4a",
  2775 => x"c2",
  2776 => x"92",
  2777 => x"c1",
  2778 => x"c3",
  2779 => x"ca",
  2780 => x"82",
  2781 => x"9f",
  2782 => x"6a",
  2783 => x"49",
  2784 => x"eb",
  2785 => x"fc",
  2786 => x"87",
  2787 => x"70",
  2788 => x"4d",
  2789 => x"75",
  2790 => x"48",
  2791 => x"ed",
  2792 => x"c9",
  2793 => x"87",
  2794 => x"0e",
  2795 => x"5e",
  2796 => x"5b",
  2797 => x"5c",
  2798 => x"5d",
  2799 => x"0e",
  2800 => x"f4",
  2801 => x"86",
  2802 => x"71",
  2803 => x"4c",
  2804 => x"c0",
  2805 => x"4b",
  2806 => x"c1",
  2807 => x"cc",
  2808 => x"c2",
  2809 => x"48",
  2810 => x"ff",
  2811 => x"78",
  2812 => x"c1",
  2813 => x"cb",
  2814 => x"e6",
  2815 => x"bf",
  2816 => x"4d",
  2817 => x"c1",
  2818 => x"cb",
  2819 => x"ea",
  2820 => x"bf",
  2821 => x"7e",
  2822 => x"c1",
  2823 => x"cb",
  2824 => x"d2",
  2825 => x"bf",
  2826 => x"02",
  2827 => x"c9",
  2828 => x"87",
  2829 => x"c1",
  2830 => x"cb",
  2831 => x"ca",
  2832 => x"bf",
  2833 => x"4a",
  2834 => x"c4",
  2835 => x"32",
  2836 => x"c7",
  2837 => x"87",
  2838 => x"c1",
  2839 => x"cb",
  2840 => x"ee",
  2841 => x"bf",
  2842 => x"4a",
  2843 => x"c4",
  2844 => x"32",
  2845 => x"c8",
  2846 => x"a6",
  2847 => x"5a",
  2848 => x"c8",
  2849 => x"a6",
  2850 => x"48",
  2851 => x"c0",
  2852 => x"78",
  2853 => x"c4",
  2854 => x"66",
  2855 => x"48",
  2856 => x"c0",
  2857 => x"a8",
  2858 => x"06",
  2859 => x"c3",
  2860 => x"cf",
  2861 => x"87",
  2862 => x"c8",
  2863 => x"66",
  2864 => x"49",
  2865 => x"cf",
  2866 => x"99",
  2867 => x"05",
  2868 => x"c0",
  2869 => x"e3",
  2870 => x"87",
  2871 => x"6e",
  2872 => x"1e",
  2873 => x"c0",
  2874 => x"e8",
  2875 => x"d5",
  2876 => x"1e",
  2877 => x"d4",
  2878 => x"c7",
  2879 => x"87",
  2880 => x"c1",
  2881 => x"c3",
  2882 => x"ca",
  2883 => x"1e",
  2884 => x"cc",
  2885 => x"66",
  2886 => x"49",
  2887 => x"48",
  2888 => x"c1",
  2889 => x"80",
  2890 => x"d0",
  2891 => x"a6",
  2892 => x"58",
  2893 => x"71",
  2894 => x"49",
  2895 => x"e7",
  2896 => x"c5",
  2897 => x"87",
  2898 => x"cc",
  2899 => x"86",
  2900 => x"c1",
  2901 => x"c3",
  2902 => x"ca",
  2903 => x"4b",
  2904 => x"c3",
  2905 => x"87",
  2906 => x"c0",
  2907 => x"e0",
  2908 => x"83",
  2909 => x"97",
  2910 => x"6b",
  2911 => x"49",
  2912 => x"71",
  2913 => x"99",
  2914 => x"02",
  2915 => x"c2",
  2916 => x"c5",
  2917 => x"87",
  2918 => x"97",
  2919 => x"6b",
  2920 => x"49",
  2921 => x"c3",
  2922 => x"e5",
  2923 => x"a9",
  2924 => x"02",
  2925 => x"c1",
  2926 => x"fb",
  2927 => x"87",
  2928 => x"cb",
  2929 => x"a3",
  2930 => x"49",
  2931 => x"97",
  2932 => x"69",
  2933 => x"49",
  2934 => x"d8",
  2935 => x"99",
  2936 => x"05",
  2937 => x"c1",
  2938 => x"ef",
  2939 => x"87",
  2940 => x"cb",
  2941 => x"1e",
  2942 => x"c0",
  2943 => x"e0",
  2944 => x"66",
  2945 => x"1e",
  2946 => x"73",
  2947 => x"49",
  2948 => x"e9",
  2949 => x"f2",
  2950 => x"87",
  2951 => x"c8",
  2952 => x"86",
  2953 => x"70",
  2954 => x"98",
  2955 => x"05",
  2956 => x"c1",
  2957 => x"dc",
  2958 => x"87",
  2959 => x"dc",
  2960 => x"a3",
  2961 => x"4a",
  2962 => x"6a",
  2963 => x"49",
  2964 => x"e8",
  2965 => x"ce",
  2966 => x"87",
  2967 => x"70",
  2968 => x"4a",
  2969 => x"c4",
  2970 => x"a4",
  2971 => x"49",
  2972 => x"72",
  2973 => x"79",
  2974 => x"da",
  2975 => x"a3",
  2976 => x"4a",
  2977 => x"9f",
  2978 => x"6a",
  2979 => x"49",
  2980 => x"e8",
  2981 => x"f8",
  2982 => x"87",
  2983 => x"c4",
  2984 => x"a6",
  2985 => x"58",
  2986 => x"c1",
  2987 => x"cb",
  2988 => x"d2",
  2989 => x"bf",
  2990 => x"02",
  2991 => x"d8",
  2992 => x"87",
  2993 => x"d4",
  2994 => x"a3",
  2995 => x"4a",
  2996 => x"9f",
  2997 => x"6a",
  2998 => x"49",
  2999 => x"e8",
  3000 => x"e5",
  3001 => x"87",
  3002 => x"70",
  3003 => x"49",
  3004 => x"c0",
  3005 => x"ff",
  3006 => x"ff",
  3007 => x"99",
  3008 => x"71",
  3009 => x"48",
  3010 => x"d0",
  3011 => x"30",
  3012 => x"c8",
  3013 => x"a6",
  3014 => x"58",
  3015 => x"c5",
  3016 => x"87",
  3017 => x"c4",
  3018 => x"a6",
  3019 => x"48",
  3020 => x"c0",
  3021 => x"78",
  3022 => x"c4",
  3023 => x"66",
  3024 => x"4a",
  3025 => x"6e",
  3026 => x"82",
  3027 => x"c8",
  3028 => x"a4",
  3029 => x"49",
  3030 => x"72",
  3031 => x"79",
  3032 => x"c0",
  3033 => x"7c",
  3034 => x"dc",
  3035 => x"66",
  3036 => x"1e",
  3037 => x"c0",
  3038 => x"e8",
  3039 => x"f2",
  3040 => x"1e",
  3041 => x"d1",
  3042 => x"e3",
  3043 => x"87",
  3044 => x"c8",
  3045 => x"86",
  3046 => x"c1",
  3047 => x"48",
  3048 => x"c1",
  3049 => x"d0",
  3050 => x"87",
  3051 => x"c8",
  3052 => x"66",
  3053 => x"48",
  3054 => x"c1",
  3055 => x"80",
  3056 => x"cc",
  3057 => x"a6",
  3058 => x"58",
  3059 => x"c8",
  3060 => x"66",
  3061 => x"48",
  3062 => x"c4",
  3063 => x"66",
  3064 => x"a8",
  3065 => x"04",
  3066 => x"fc",
  3067 => x"f1",
  3068 => x"87",
  3069 => x"c1",
  3070 => x"cb",
  3071 => x"d2",
  3072 => x"bf",
  3073 => x"02",
  3074 => x"c0",
  3075 => x"f4",
  3076 => x"87",
  3077 => x"75",
  3078 => x"49",
  3079 => x"f9",
  3080 => x"e0",
  3081 => x"87",
  3082 => x"70",
  3083 => x"4d",
  3084 => x"75",
  3085 => x"1e",
  3086 => x"c0",
  3087 => x"e9",
  3088 => x"c3",
  3089 => x"1e",
  3090 => x"d0",
  3091 => x"f2",
  3092 => x"87",
  3093 => x"c8",
  3094 => x"86",
  3095 => x"75",
  3096 => x"49",
  3097 => x"cf",
  3098 => x"ff",
  3099 => x"ff",
  3100 => x"ff",
  3101 => x"f8",
  3102 => x"99",
  3103 => x"a9",
  3104 => x"02",
  3105 => x"d6",
  3106 => x"87",
  3107 => x"75",
  3108 => x"49",
  3109 => x"c2",
  3110 => x"89",
  3111 => x"c1",
  3112 => x"cb",
  3113 => x"ca",
  3114 => x"bf",
  3115 => x"91",
  3116 => x"c1",
  3117 => x"cb",
  3118 => x"e2",
  3119 => x"bf",
  3120 => x"48",
  3121 => x"71",
  3122 => x"80",
  3123 => x"c4",
  3124 => x"a6",
  3125 => x"58",
  3126 => x"fb",
  3127 => x"e7",
  3128 => x"87",
  3129 => x"c0",
  3130 => x"48",
  3131 => x"f4",
  3132 => x"8e",
  3133 => x"e7",
  3134 => x"f3",
  3135 => x"87",
  3136 => x"0e",
  3137 => x"5e",
  3138 => x"5b",
  3139 => x"5c",
  3140 => x"5d",
  3141 => x"0e",
  3142 => x"1e",
  3143 => x"71",
  3144 => x"4b",
  3145 => x"73",
  3146 => x"1e",
  3147 => x"c1",
  3148 => x"cc",
  3149 => x"c6",
  3150 => x"49",
  3151 => x"fa",
  3152 => x"d8",
  3153 => x"87",
  3154 => x"c4",
  3155 => x"86",
  3156 => x"70",
  3157 => x"98",
  3158 => x"02",
  3159 => x"c1",
  3160 => x"f7",
  3161 => x"87",
  3162 => x"c1",
  3163 => x"cc",
  3164 => x"ca",
  3165 => x"bf",
  3166 => x"49",
  3167 => x"c7",
  3168 => x"ff",
  3169 => x"81",
  3170 => x"c9",
  3171 => x"29",
  3172 => x"c4",
  3173 => x"a6",
  3174 => x"59",
  3175 => x"c0",
  3176 => x"4d",
  3177 => x"4c",
  3178 => x"6e",
  3179 => x"48",
  3180 => x"c0",
  3181 => x"b7",
  3182 => x"a8",
  3183 => x"06",
  3184 => x"c1",
  3185 => x"ed",
  3186 => x"87",
  3187 => x"c1",
  3188 => x"cb",
  3189 => x"e2",
  3190 => x"bf",
  3191 => x"49",
  3192 => x"c1",
  3193 => x"cc",
  3194 => x"ce",
  3195 => x"bf",
  3196 => x"4a",
  3197 => x"c2",
  3198 => x"8a",
  3199 => x"c1",
  3200 => x"cb",
  3201 => x"ca",
  3202 => x"bf",
  3203 => x"92",
  3204 => x"72",
  3205 => x"a1",
  3206 => x"49",
  3207 => x"c1",
  3208 => x"cb",
  3209 => x"ce",
  3210 => x"bf",
  3211 => x"4a",
  3212 => x"74",
  3213 => x"9a",
  3214 => x"72",
  3215 => x"a1",
  3216 => x"49",
  3217 => x"d4",
  3218 => x"66",
  3219 => x"1e",
  3220 => x"71",
  3221 => x"49",
  3222 => x"e1",
  3223 => x"fe",
  3224 => x"87",
  3225 => x"c4",
  3226 => x"86",
  3227 => x"70",
  3228 => x"98",
  3229 => x"05",
  3230 => x"c5",
  3231 => x"87",
  3232 => x"c0",
  3233 => x"48",
  3234 => x"c1",
  3235 => x"c0",
  3236 => x"87",
  3237 => x"c1",
  3238 => x"84",
  3239 => x"c1",
  3240 => x"cb",
  3241 => x"ce",
  3242 => x"bf",
  3243 => x"49",
  3244 => x"74",
  3245 => x"99",
  3246 => x"05",
  3247 => x"cc",
  3248 => x"87",
  3249 => x"c1",
  3250 => x"cc",
  3251 => x"ce",
  3252 => x"bf",
  3253 => x"49",
  3254 => x"f6",
  3255 => x"f1",
  3256 => x"87",
  3257 => x"c1",
  3258 => x"cc",
  3259 => x"d2",
  3260 => x"58",
  3261 => x"d4",
  3262 => x"66",
  3263 => x"48",
  3264 => x"c8",
  3265 => x"c0",
  3266 => x"80",
  3267 => x"d8",
  3268 => x"a6",
  3269 => x"58",
  3270 => x"c1",
  3271 => x"85",
  3272 => x"6e",
  3273 => x"b7",
  3274 => x"ad",
  3275 => x"04",
  3276 => x"fe",
  3277 => x"e4",
  3278 => x"87",
  3279 => x"cf",
  3280 => x"87",
  3281 => x"73",
  3282 => x"1e",
  3283 => x"c0",
  3284 => x"e9",
  3285 => x"db",
  3286 => x"1e",
  3287 => x"cd",
  3288 => x"ed",
  3289 => x"87",
  3290 => x"c8",
  3291 => x"86",
  3292 => x"c0",
  3293 => x"48",
  3294 => x"c5",
  3295 => x"87",
  3296 => x"c1",
  3297 => x"cc",
  3298 => x"ca",
  3299 => x"bf",
  3300 => x"48",
  3301 => x"26",
  3302 => x"e5",
  3303 => x"ca",
  3304 => x"87",
  3305 => x"1e",
  3306 => x"c0",
  3307 => x"f6",
  3308 => x"e8",
  3309 => x"c0",
  3310 => x"c0",
  3311 => x"09",
  3312 => x"97",
  3313 => x"79",
  3314 => x"09",
  3315 => x"71",
  3316 => x"48",
  3317 => x"26",
  3318 => x"4f",
  3319 => x"0e",
  3320 => x"5e",
  3321 => x"5b",
  3322 => x"5c",
  3323 => x"0e",
  3324 => x"71",
  3325 => x"4b",
  3326 => x"c0",
  3327 => x"4c",
  3328 => x"13",
  3329 => x"4a",
  3330 => x"72",
  3331 => x"9a",
  3332 => x"02",
  3333 => x"ce",
  3334 => x"87",
  3335 => x"72",
  3336 => x"49",
  3337 => x"ff",
  3338 => x"dd",
  3339 => x"87",
  3340 => x"c1",
  3341 => x"84",
  3342 => x"13",
  3343 => x"4a",
  3344 => x"72",
  3345 => x"9a",
  3346 => x"05",
  3347 => x"f2",
  3348 => x"87",
  3349 => x"74",
  3350 => x"48",
  3351 => x"c2",
  3352 => x"87",
  3353 => x"26",
  3354 => x"4d",
  3355 => x"26",
  3356 => x"4c",
  3357 => x"26",
  3358 => x"4b",
  3359 => x"26",
  3360 => x"4f",
  3361 => x"0e",
  3362 => x"5e",
  3363 => x"5b",
  3364 => x"5c",
  3365 => x"5d",
  3366 => x"0e",
  3367 => x"71",
  3368 => x"4b",
  3369 => x"73",
  3370 => x"4c",
  3371 => x"d0",
  3372 => x"66",
  3373 => x"48",
  3374 => x"c2",
  3375 => x"28",
  3376 => x"d4",
  3377 => x"a6",
  3378 => x"58",
  3379 => x"d0",
  3380 => x"66",
  3381 => x"49",
  3382 => x"48",
  3383 => x"c1",
  3384 => x"88",
  3385 => x"d4",
  3386 => x"a6",
  3387 => x"58",
  3388 => x"71",
  3389 => x"99",
  3390 => x"02",
  3391 => x"c1",
  3392 => x"c4",
  3393 => x"87",
  3394 => x"24",
  3395 => x"4d",
  3396 => x"c0",
  3397 => x"4b",
  3398 => x"75",
  3399 => x"4a",
  3400 => x"dc",
  3401 => x"2a",
  3402 => x"c0",
  3403 => x"f0",
  3404 => x"82",
  3405 => x"c0",
  3406 => x"f9",
  3407 => x"aa",
  3408 => x"06",
  3409 => x"c2",
  3410 => x"87",
  3411 => x"c7",
  3412 => x"82",
  3413 => x"72",
  3414 => x"49",
  3415 => x"fe",
  3416 => x"cf",
  3417 => x"87",
  3418 => x"c4",
  3419 => x"35",
  3420 => x"c1",
  3421 => x"83",
  3422 => x"c8",
  3423 => x"b7",
  3424 => x"ab",
  3425 => x"04",
  3426 => x"e2",
  3427 => x"87",
  3428 => x"c0",
  3429 => x"e0",
  3430 => x"49",
  3431 => x"fd",
  3432 => x"ff",
  3433 => x"87",
  3434 => x"d0",
  3435 => x"66",
  3436 => x"49",
  3437 => x"c3",
  3438 => x"99",
  3439 => x"05",
  3440 => x"c5",
  3441 => x"87",
  3442 => x"ca",
  3443 => x"49",
  3444 => x"fd",
  3445 => x"f2",
  3446 => x"87",
  3447 => x"d0",
  3448 => x"66",
  3449 => x"49",
  3450 => x"48",
  3451 => x"c1",
  3452 => x"88",
  3453 => x"d4",
  3454 => x"a6",
  3455 => x"58",
  3456 => x"71",
  3457 => x"99",
  3458 => x"05",
  3459 => x"fe",
  3460 => x"fc",
  3461 => x"87",
  3462 => x"ca",
  3463 => x"49",
  3464 => x"fd",
  3465 => x"de",
  3466 => x"87",
  3467 => x"26",
  3468 => x"4d",
  3469 => x"26",
  3470 => x"4c",
  3471 => x"26",
  3472 => x"4b",
  3473 => x"26",
  3474 => x"4f",
  3475 => x"0e",
  3476 => x"5e",
  3477 => x"5b",
  3478 => x"5c",
  3479 => x"5d",
  3480 => x"0e",
  3481 => x"fc",
  3482 => x"86",
  3483 => x"71",
  3484 => x"4a",
  3485 => x"c0",
  3486 => x"e0",
  3487 => x"66",
  3488 => x"4c",
  3489 => x"c1",
  3490 => x"cc",
  3491 => x"d2",
  3492 => x"4b",
  3493 => x"c0",
  3494 => x"7e",
  3495 => x"72",
  3496 => x"9a",
  3497 => x"05",
  3498 => x"ce",
  3499 => x"87",
  3500 => x"c1",
  3501 => x"cc",
  3502 => x"d3",
  3503 => x"4b",
  3504 => x"c1",
  3505 => x"cc",
  3506 => x"d2",
  3507 => x"48",
  3508 => x"c0",
  3509 => x"f0",
  3510 => x"50",
  3511 => x"c1",
  3512 => x"d2",
  3513 => x"87",
  3514 => x"72",
  3515 => x"9a",
  3516 => x"02",
  3517 => x"c0",
  3518 => x"e9",
  3519 => x"87",
  3520 => x"d4",
  3521 => x"66",
  3522 => x"4d",
  3523 => x"72",
  3524 => x"1e",
  3525 => x"72",
  3526 => x"49",
  3527 => x"75",
  3528 => x"4a",
  3529 => x"ca",
  3530 => x"cf",
  3531 => x"87",
  3532 => x"26",
  3533 => x"4a",
  3534 => x"c0",
  3535 => x"f8",
  3536 => x"fd",
  3537 => x"81",
  3538 => x"11",
  3539 => x"53",
  3540 => x"71",
  3541 => x"1e",
  3542 => x"72",
  3543 => x"49",
  3544 => x"75",
  3545 => x"4a",
  3546 => x"c9",
  3547 => x"fe",
  3548 => x"87",
  3549 => x"70",
  3550 => x"4a",
  3551 => x"26",
  3552 => x"49",
  3553 => x"c1",
  3554 => x"8c",
  3555 => x"72",
  3556 => x"9a",
  3557 => x"05",
  3558 => x"ff",
  3559 => x"da",
  3560 => x"87",
  3561 => x"c0",
  3562 => x"b7",
  3563 => x"ac",
  3564 => x"06",
  3565 => x"dd",
  3566 => x"87",
  3567 => x"c0",
  3568 => x"e4",
  3569 => x"66",
  3570 => x"02",
  3571 => x"c5",
  3572 => x"87",
  3573 => x"c0",
  3574 => x"f0",
  3575 => x"4a",
  3576 => x"c3",
  3577 => x"87",
  3578 => x"c0",
  3579 => x"e0",
  3580 => x"4a",
  3581 => x"73",
  3582 => x"0a",
  3583 => x"97",
  3584 => x"7a",
  3585 => x"0a",
  3586 => x"c1",
  3587 => x"83",
  3588 => x"8c",
  3589 => x"c0",
  3590 => x"b7",
  3591 => x"ac",
  3592 => x"01",
  3593 => x"ff",
  3594 => x"e3",
  3595 => x"87",
  3596 => x"c1",
  3597 => x"cc",
  3598 => x"d2",
  3599 => x"ab",
  3600 => x"02",
  3601 => x"de",
  3602 => x"87",
  3603 => x"d8",
  3604 => x"66",
  3605 => x"4c",
  3606 => x"dc",
  3607 => x"66",
  3608 => x"1e",
  3609 => x"c1",
  3610 => x"8b",
  3611 => x"97",
  3612 => x"6b",
  3613 => x"49",
  3614 => x"74",
  3615 => x"0f",
  3616 => x"c4",
  3617 => x"86",
  3618 => x"6e",
  3619 => x"48",
  3620 => x"c1",
  3621 => x"80",
  3622 => x"c4",
  3623 => x"a6",
  3624 => x"58",
  3625 => x"c1",
  3626 => x"cc",
  3627 => x"d2",
  3628 => x"ab",
  3629 => x"05",
  3630 => x"ff",
  3631 => x"e5",
  3632 => x"87",
  3633 => x"6e",
  3634 => x"48",
  3635 => x"fc",
  3636 => x"8e",
  3637 => x"26",
  3638 => x"4d",
  3639 => x"26",
  3640 => x"4c",
  3641 => x"26",
  3642 => x"4b",
  3643 => x"26",
  3644 => x"4f",
  3645 => x"30",
  3646 => x"31",
  3647 => x"32",
  3648 => x"33",
  3649 => x"34",
  3650 => x"35",
  3651 => x"36",
  3652 => x"37",
  3653 => x"38",
  3654 => x"39",
  3655 => x"41",
  3656 => x"42",
  3657 => x"43",
  3658 => x"44",
  3659 => x"45",
  3660 => x"46",
  3661 => x"00",
  3662 => x"0e",
  3663 => x"5e",
  3664 => x"5b",
  3665 => x"5c",
  3666 => x"5d",
  3667 => x"0e",
  3668 => x"71",
  3669 => x"4b",
  3670 => x"ff",
  3671 => x"4d",
  3672 => x"13",
  3673 => x"4c",
  3674 => x"74",
  3675 => x"9c",
  3676 => x"02",
  3677 => x"d8",
  3678 => x"87",
  3679 => x"c1",
  3680 => x"85",
  3681 => x"d4",
  3682 => x"66",
  3683 => x"1e",
  3684 => x"74",
  3685 => x"49",
  3686 => x"d4",
  3687 => x"66",
  3688 => x"0f",
  3689 => x"c4",
  3690 => x"86",
  3691 => x"74",
  3692 => x"a8",
  3693 => x"05",
  3694 => x"c7",
  3695 => x"87",
  3696 => x"13",
  3697 => x"4c",
  3698 => x"74",
  3699 => x"9c",
  3700 => x"05",
  3701 => x"e8",
  3702 => x"87",
  3703 => x"75",
  3704 => x"48",
  3705 => x"26",
  3706 => x"4d",
  3707 => x"26",
  3708 => x"4c",
  3709 => x"26",
  3710 => x"4b",
  3711 => x"26",
  3712 => x"4f",
  3713 => x"0e",
  3714 => x"5e",
  3715 => x"5b",
  3716 => x"5c",
  3717 => x"5d",
  3718 => x"0e",
  3719 => x"e8",
  3720 => x"86",
  3721 => x"c4",
  3722 => x"a6",
  3723 => x"59",
  3724 => x"c0",
  3725 => x"e8",
  3726 => x"66",
  3727 => x"4d",
  3728 => x"c0",
  3729 => x"4c",
  3730 => x"c8",
  3731 => x"a6",
  3732 => x"48",
  3733 => x"c0",
  3734 => x"78",
  3735 => x"6e",
  3736 => x"97",
  3737 => x"bf",
  3738 => x"4b",
  3739 => x"6e",
  3740 => x"48",
  3741 => x"c1",
  3742 => x"80",
  3743 => x"c4",
  3744 => x"a6",
  3745 => x"58",
  3746 => x"73",
  3747 => x"9b",
  3748 => x"02",
  3749 => x"c6",
  3750 => x"d3",
  3751 => x"87",
  3752 => x"c8",
  3753 => x"66",
  3754 => x"02",
  3755 => x"c5",
  3756 => x"db",
  3757 => x"87",
  3758 => x"cc",
  3759 => x"a6",
  3760 => x"48",
  3761 => x"c0",
  3762 => x"78",
  3763 => x"fc",
  3764 => x"80",
  3765 => x"c0",
  3766 => x"78",
  3767 => x"73",
  3768 => x"4a",
  3769 => x"c0",
  3770 => x"e0",
  3771 => x"8a",
  3772 => x"02",
  3773 => x"c3",
  3774 => x"c6",
  3775 => x"87",
  3776 => x"c3",
  3777 => x"8a",
  3778 => x"02",
  3779 => x"c3",
  3780 => x"c0",
  3781 => x"87",
  3782 => x"c2",
  3783 => x"8a",
  3784 => x"02",
  3785 => x"c2",
  3786 => x"e8",
  3787 => x"87",
  3788 => x"c2",
  3789 => x"8a",
  3790 => x"02",
  3791 => x"c2",
  3792 => x"f4",
  3793 => x"87",
  3794 => x"c4",
  3795 => x"8a",
  3796 => x"02",
  3797 => x"c2",
  3798 => x"ee",
  3799 => x"87",
  3800 => x"c2",
  3801 => x"8a",
  3802 => x"02",
  3803 => x"c2",
  3804 => x"e8",
  3805 => x"87",
  3806 => x"c3",
  3807 => x"8a",
  3808 => x"02",
  3809 => x"c2",
  3810 => x"ea",
  3811 => x"87",
  3812 => x"d4",
  3813 => x"8a",
  3814 => x"02",
  3815 => x"c0",
  3816 => x"f6",
  3817 => x"87",
  3818 => x"d4",
  3819 => x"8a",
  3820 => x"02",
  3821 => x"c1",
  3822 => x"c0",
  3823 => x"87",
  3824 => x"ca",
  3825 => x"8a",
  3826 => x"02",
  3827 => x"c0",
  3828 => x"f2",
  3829 => x"87",
  3830 => x"c1",
  3831 => x"8a",
  3832 => x"02",
  3833 => x"c1",
  3834 => x"e1",
  3835 => x"87",
  3836 => x"c1",
  3837 => x"8a",
  3838 => x"02",
  3839 => x"df",
  3840 => x"87",
  3841 => x"c8",
  3842 => x"8a",
  3843 => x"02",
  3844 => x"c1",
  3845 => x"ce",
  3846 => x"87",
  3847 => x"c4",
  3848 => x"8a",
  3849 => x"02",
  3850 => x"c0",
  3851 => x"e3",
  3852 => x"87",
  3853 => x"c3",
  3854 => x"8a",
  3855 => x"02",
  3856 => x"c0",
  3857 => x"e5",
  3858 => x"87",
  3859 => x"c2",
  3860 => x"8a",
  3861 => x"02",
  3862 => x"c8",
  3863 => x"87",
  3864 => x"c3",
  3865 => x"8a",
  3866 => x"02",
  3867 => x"d3",
  3868 => x"87",
  3869 => x"c1",
  3870 => x"fa",
  3871 => x"87",
  3872 => x"cc",
  3873 => x"a6",
  3874 => x"48",
  3875 => x"ca",
  3876 => x"78",
  3877 => x"c2",
  3878 => x"d2",
  3879 => x"87",
  3880 => x"cc",
  3881 => x"a6",
  3882 => x"48",
  3883 => x"c2",
  3884 => x"78",
  3885 => x"c2",
  3886 => x"ca",
  3887 => x"87",
  3888 => x"cc",
  3889 => x"a6",
  3890 => x"48",
  3891 => x"d0",
  3892 => x"78",
  3893 => x"c2",
  3894 => x"c2",
  3895 => x"87",
  3896 => x"c0",
  3897 => x"f0",
  3898 => x"66",
  3899 => x"1e",
  3900 => x"c0",
  3901 => x"f0",
  3902 => x"66",
  3903 => x"1e",
  3904 => x"c4",
  3905 => x"85",
  3906 => x"75",
  3907 => x"4a",
  3908 => x"c4",
  3909 => x"8a",
  3910 => x"6a",
  3911 => x"49",
  3912 => x"fc",
  3913 => x"c3",
  3914 => x"87",
  3915 => x"c8",
  3916 => x"86",
  3917 => x"70",
  3918 => x"49",
  3919 => x"71",
  3920 => x"a4",
  3921 => x"4c",
  3922 => x"c1",
  3923 => x"e5",
  3924 => x"87",
  3925 => x"c8",
  3926 => x"a6",
  3927 => x"48",
  3928 => x"c1",
  3929 => x"78",
  3930 => x"c1",
  3931 => x"dd",
  3932 => x"87",
  3933 => x"c0",
  3934 => x"f0",
  3935 => x"66",
  3936 => x"1e",
  3937 => x"c4",
  3938 => x"85",
  3939 => x"75",
  3940 => x"4a",
  3941 => x"c4",
  3942 => x"8a",
  3943 => x"6a",
  3944 => x"49",
  3945 => x"c0",
  3946 => x"f0",
  3947 => x"66",
  3948 => x"0f",
  3949 => x"c4",
  3950 => x"86",
  3951 => x"c1",
  3952 => x"84",
  3953 => x"c1",
  3954 => x"c6",
  3955 => x"87",
  3956 => x"c0",
  3957 => x"f0",
  3958 => x"66",
  3959 => x"1e",
  3960 => x"c0",
  3961 => x"e5",
  3962 => x"49",
  3963 => x"c0",
  3964 => x"f0",
  3965 => x"66",
  3966 => x"0f",
  3967 => x"c4",
  3968 => x"86",
  3969 => x"c1",
  3970 => x"84",
  3971 => x"c0",
  3972 => x"f4",
  3973 => x"87",
  3974 => x"c8",
  3975 => x"a6",
  3976 => x"48",
  3977 => x"c1",
  3978 => x"78",
  3979 => x"c0",
  3980 => x"ec",
  3981 => x"87",
  3982 => x"d0",
  3983 => x"a6",
  3984 => x"48",
  3985 => x"c1",
  3986 => x"78",
  3987 => x"f8",
  3988 => x"80",
  3989 => x"c1",
  3990 => x"78",
  3991 => x"c0",
  3992 => x"e0",
  3993 => x"87",
  3994 => x"c0",
  3995 => x"f0",
  3996 => x"ab",
  3997 => x"06",
  3998 => x"da",
  3999 => x"87",
  4000 => x"c0",
  4001 => x"f9",
  4002 => x"ab",
  4003 => x"03",
  4004 => x"d4",
  4005 => x"87",
  4006 => x"d4",
  4007 => x"66",
  4008 => x"49",
  4009 => x"ca",
  4010 => x"91",
  4011 => x"73",
  4012 => x"4a",
  4013 => x"c0",
  4014 => x"f0",
  4015 => x"8a",
  4016 => x"d4",
  4017 => x"a6",
  4018 => x"48",
  4019 => x"72",
  4020 => x"a1",
  4021 => x"78",
  4022 => x"f4",
  4023 => x"80",
  4024 => x"c1",
  4025 => x"78",
  4026 => x"cc",
  4027 => x"66",
  4028 => x"02",
  4029 => x"c1",
  4030 => x"ea",
  4031 => x"87",
  4032 => x"c4",
  4033 => x"85",
  4034 => x"75",
  4035 => x"49",
  4036 => x"c4",
  4037 => x"89",
  4038 => x"a6",
  4039 => x"48",
  4040 => x"69",
  4041 => x"78",
  4042 => x"c1",
  4043 => x"e4",
  4044 => x"ab",
  4045 => x"05",
  4046 => x"d8",
  4047 => x"87",
  4048 => x"c4",
  4049 => x"66",
  4050 => x"48",
  4051 => x"c0",
  4052 => x"b7",
  4053 => x"a8",
  4054 => x"03",
  4055 => x"cf",
  4056 => x"87",
  4057 => x"c0",
  4058 => x"ed",
  4059 => x"49",
  4060 => x"f4",
  4061 => x"ca",
  4062 => x"87",
  4063 => x"c4",
  4064 => x"66",
  4065 => x"48",
  4066 => x"c0",
  4067 => x"08",
  4068 => x"88",
  4069 => x"c8",
  4070 => x"a6",
  4071 => x"58",
  4072 => x"d0",
  4073 => x"66",
  4074 => x"1e",
  4075 => x"d8",
  4076 => x"66",
  4077 => x"1e",
  4078 => x"c0",
  4079 => x"f8",
  4080 => x"66",
  4081 => x"1e",
  4082 => x"c0",
  4083 => x"f8",
  4084 => x"66",
  4085 => x"1e",
  4086 => x"dc",
  4087 => x"66",
  4088 => x"1e",
  4089 => x"d8",
  4090 => x"66",
  4091 => x"49",
  4092 => x"f6",
  4093 => x"d4",
  4094 => x"87",
  4095 => x"d4",
  4096 => x"86",
  4097 => x"70",
  4098 => x"49",
  4099 => x"71",
  4100 => x"a4",
  4101 => x"4c",
  4102 => x"c0",
  4103 => x"e1",
  4104 => x"87",
  4105 => x"c0",
  4106 => x"e5",
  4107 => x"ab",
  4108 => x"05",
  4109 => x"cf",
  4110 => x"87",
  4111 => x"d0",
  4112 => x"a6",
  4113 => x"48",
  4114 => x"c0",
  4115 => x"78",
  4116 => x"c4",
  4117 => x"80",
  4118 => x"c0",
  4119 => x"78",
  4120 => x"f4",
  4121 => x"80",
  4122 => x"c1",
  4123 => x"78",
  4124 => x"cc",
  4125 => x"87",
  4126 => x"c0",
  4127 => x"f0",
  4128 => x"66",
  4129 => x"1e",
  4130 => x"73",
  4131 => x"49",
  4132 => x"c0",
  4133 => x"f0",
  4134 => x"66",
  4135 => x"0f",
  4136 => x"c4",
  4137 => x"86",
  4138 => x"6e",
  4139 => x"97",
  4140 => x"bf",
  4141 => x"4b",
  4142 => x"6e",
  4143 => x"48",
  4144 => x"c1",
  4145 => x"80",
  4146 => x"c4",
  4147 => x"a6",
  4148 => x"58",
  4149 => x"73",
  4150 => x"9b",
  4151 => x"05",
  4152 => x"f9",
  4153 => x"ed",
  4154 => x"87",
  4155 => x"74",
  4156 => x"48",
  4157 => x"e8",
  4158 => x"8e",
  4159 => x"26",
  4160 => x"4d",
  4161 => x"26",
  4162 => x"4c",
  4163 => x"26",
  4164 => x"4b",
  4165 => x"26",
  4166 => x"4f",
  4167 => x"1e",
  4168 => x"c0",
  4169 => x"1e",
  4170 => x"c0",
  4171 => x"f3",
  4172 => x"e9",
  4173 => x"1e",
  4174 => x"d0",
  4175 => x"a6",
  4176 => x"1e",
  4177 => x"d0",
  4178 => x"66",
  4179 => x"49",
  4180 => x"f8",
  4181 => x"ea",
  4182 => x"87",
  4183 => x"f4",
  4184 => x"8e",
  4185 => x"26",
  4186 => x"4f",
  4187 => x"1e",
  4188 => x"73",
  4189 => x"1e",
  4190 => x"72",
  4191 => x"9a",
  4192 => x"02",
  4193 => x"c0",
  4194 => x"e7",
  4195 => x"87",
  4196 => x"c0",
  4197 => x"48",
  4198 => x"c1",
  4199 => x"4b",
  4200 => x"72",
  4201 => x"a9",
  4202 => x"06",
  4203 => x"d1",
  4204 => x"87",
  4205 => x"72",
  4206 => x"82",
  4207 => x"06",
  4208 => x"c9",
  4209 => x"87",
  4210 => x"73",
  4211 => x"83",
  4212 => x"72",
  4213 => x"a9",
  4214 => x"01",
  4215 => x"f4",
  4216 => x"87",
  4217 => x"c3",
  4218 => x"87",
  4219 => x"c1",
  4220 => x"b2",
  4221 => x"3a",
  4222 => x"72",
  4223 => x"a9",
  4224 => x"03",
  4225 => x"89",
  4226 => x"73",
  4227 => x"80",
  4228 => x"07",
  4229 => x"c1",
  4230 => x"2a",
  4231 => x"2b",
  4232 => x"05",
  4233 => x"f3",
  4234 => x"87",
  4235 => x"26",
  4236 => x"4b",
  4237 => x"26",
  4238 => x"4f",
  4239 => x"1e",
  4240 => x"75",
  4241 => x"1e",
  4242 => x"c4",
  4243 => x"4d",
  4244 => x"71",
  4245 => x"b7",
  4246 => x"a1",
  4247 => x"04",
  4248 => x"ff",
  4249 => x"b9",
  4250 => x"c1",
  4251 => x"81",
  4252 => x"c3",
  4253 => x"bd",
  4254 => x"07",
  4255 => x"72",
  4256 => x"b7",
  4257 => x"a2",
  4258 => x"04",
  4259 => x"ff",
  4260 => x"ba",
  4261 => x"c1",
  4262 => x"82",
  4263 => x"c1",
  4264 => x"bd",
  4265 => x"07",
  4266 => x"fe",
  4267 => x"ee",
  4268 => x"87",
  4269 => x"c1",
  4270 => x"2d",
  4271 => x"04",
  4272 => x"ff",
  4273 => x"b8",
  4274 => x"c1",
  4275 => x"80",
  4276 => x"07",
  4277 => x"2d",
  4278 => x"04",
  4279 => x"ff",
  4280 => x"b9",
  4281 => x"c1",
  4282 => x"81",
  4283 => x"07",
  4284 => x"26",
  4285 => x"4d",
  4286 => x"26",
  4287 => x"4f",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;

