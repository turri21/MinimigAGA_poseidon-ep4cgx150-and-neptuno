library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM-2 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111";
	-- Second port
	addr2 : in std_logic_vector(maxAddrBitBRAM-2 downto 0) := (others=>'0');
	q2 : out std_logic_vector(31 downto 0);
	d2 : in std_logic_vector(31 downto 0) := X"00000000";
	we2 : in std_logic := '0';
	bytesel2 : in std_logic_vector(3 downto 0) := "1111"	
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
type ram_type is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

signal ram : ram_type :=
(
     0 => (x"01",x"da",x"87",x"04"),
     1 => (x"dd",x"87",x"0e",x"58"),
     2 => (x"5e",x"59",x"5a",x"0e"),
     3 => (x"27",x"00",x"00",x"00"),
     4 => (x"29",x"0f",x"26",x"4a"),
     5 => (x"26",x"49",x"26",x"48"),
     6 => (x"ff",x"80",x"26",x"08"),
     7 => (x"4f",x"27",x"00",x"00"),
     8 => (x"00",x"2d",x"4f",x"27"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"4f",x"4f",x"00",x"fd"),
    11 => (x"87",x"c1",x"ca",x"c0"),
    12 => (x"4e",x"c9",x"c0",x"48"),
    13 => (x"c2",x"28",x"c1",x"d5"),
    14 => (x"ea",x"e5",x"d6",x"ea"),
    15 => (x"49",x"71",x"46",x"c1"),
    16 => (x"88",x"01",x"f9",x"87"),
    17 => (x"c1",x"ca",x"c0",x"49"),
    18 => (x"c1",x"c0",x"ec",x"48"),
    19 => (x"89",x"d0",x"89",x"03"),
    20 => (x"c0",x"40",x"40",x"40"),
    21 => (x"40",x"f6",x"87",x"d0"),
    22 => (x"81",x"05",x"c0",x"50"),
    23 => (x"c1",x"89",x"05",x"f9"),
    24 => (x"87",x"c1",x"c0",x"ea"),
    25 => (x"4d",x"c1",x"c0",x"ea"),
    26 => (x"4c",x"74",x"ad",x"02"),
    27 => (x"c4",x"87",x"24",x"0f"),
    28 => (x"f7",x"87",x"c2",x"dc"),
    29 => (x"87",x"c1",x"c0",x"ea"),
    30 => (x"4d",x"c1",x"c0",x"ea"),
    31 => (x"4c",x"74",x"ad",x"02"),
    32 => (x"c6",x"87",x"c4",x"8c"),
    33 => (x"6c",x"0f",x"f5",x"87"),
    34 => (x"00",x"98",x"fc",x"87"),
    35 => (x"0e",x"5e",x"5b",x"5c"),
    36 => (x"0e",x"c4",x"c0",x"c0"),
    37 => (x"c0",x"4b",x"c9",x"d0"),
    38 => (x"4c",x"c9",x"e2",x"bf"),
    39 => (x"4a",x"49",x"c1",x"8a"),
    40 => (x"71",x"99",x"02",x"cf"),
    41 => (x"87",x"74",x"49",x"c1"),
    42 => (x"84",x"11",x"53",x"72"),
    43 => (x"49",x"c1",x"8a",x"71"),
    44 => (x"99",x"05",x"f1",x"87"),
    45 => (x"c2",x"87",x"26",x"4d"),
    46 => (x"26",x"4c",x"26",x"4b"),
    47 => (x"26",x"4f",x"1e",x"73"),
    48 => (x"1e",x"71",x"4b",x"e7"),
    49 => (x"48",x"c0",x"e0",x"50"),
    50 => (x"e3",x"48",x"c8",x"50"),
    51 => (x"e3",x"48",x"c6",x"50"),
    52 => (x"e7",x"48",x"c0",x"e1"),
    53 => (x"50",x"73",x"4a",x"c8"),
    54 => (x"b7",x"2a",x"c4",x"c0"),
    55 => (x"c0",x"c0",x"49",x"ca"),
    56 => (x"81",x"72",x"51",x"73"),
    57 => (x"4a",x"c3",x"ff",x"9a"),
    58 => (x"c4",x"c0",x"c0",x"c0"),
    59 => (x"49",x"cb",x"81",x"72"),
    60 => (x"51",x"e7",x"48",x"c0"),
    61 => (x"e0",x"50",x"e3",x"48"),
    62 => (x"c8",x"50",x"e3",x"48"),
    63 => (x"c0",x"50",x"e7",x"48"),
    64 => (x"c0",x"e1",x"50",x"fe"),
    65 => (x"f4",x"87",x"1e",x"73"),
    66 => (x"1e",x"c2",x"c0",x"c0"),
    67 => (x"4b",x"0f",x"fe",x"e9"),
    68 => (x"87",x"1e",x"73",x"1e"),
    69 => (x"eb",x"48",x"c3",x"ef"),
    70 => (x"50",x"e7",x"48",x"c0"),
    71 => (x"e0",x"50",x"e3",x"48"),
    72 => (x"c8",x"50",x"e3",x"48"),
    73 => (x"c6",x"50",x"e7",x"48"),
    74 => (x"c0",x"e1",x"50",x"ff"),
    75 => (x"c2",x"48",x"c1",x"9f"),
    76 => (x"78",x"e7",x"48",x"c0"),
    77 => (x"e0",x"50",x"e3",x"48"),
    78 => (x"c4",x"50",x"e3",x"48"),
    79 => (x"c2",x"50",x"e7",x"48"),
    80 => (x"c0",x"e1",x"50",x"e7"),
    81 => (x"48",x"c0",x"e0",x"50"),
    82 => (x"e3",x"48",x"c8",x"50"),
    83 => (x"e3",x"48",x"c7",x"50"),
    84 => (x"e7",x"48",x"c0",x"e1"),
    85 => (x"50",x"fc",x"f4",x"87"),
    86 => (x"c0",x"ff",x"ff",x"49"),
    87 => (x"fd",x"df",x"87",x"c0"),
    88 => (x"fc",x"c0",x"4b",x"c8"),
    89 => (x"dc",x"49",x"c0",x"f8"),
    90 => (x"f7",x"87",x"cd",x"e5"),
    91 => (x"87",x"70",x"98",x"02"),
    92 => (x"c1",x"c3",x"87",x"c0"),
    93 => (x"ff",x"f0",x"4b",x"c8"),
    94 => (x"c5",x"49",x"c0",x"f8"),
    95 => (x"e3",x"87",x"d3",x"cf"),
    96 => (x"87",x"70",x"98",x"02"),
    97 => (x"c0",x"e6",x"87",x"c3"),
    98 => (x"f0",x"4b",x"c2",x"c0"),
    99 => (x"c0",x"1e",x"c7",x"c8"),
   100 => (x"49",x"c0",x"ea",x"d2"),
   101 => (x"87",x"c4",x"86",x"70"),
   102 => (x"98",x"02",x"c8",x"87"),
   103 => (x"c3",x"ff",x"4b",x"fd"),
   104 => (x"e4",x"87",x"d9",x"87"),
   105 => (x"c7",x"d4",x"49",x"c0"),
   106 => (x"f7",x"f6",x"87",x"d0"),
   107 => (x"87",x"c7",x"e9",x"49"),
   108 => (x"c0",x"f7",x"ed",x"87"),
   109 => (x"c7",x"87",x"c8",x"f2"),
   110 => (x"49",x"c0",x"f7",x"e4"),
   111 => (x"87",x"73",x"49",x"fb"),
   112 => (x"fc",x"87",x"fe",x"da"),
   113 => (x"87",x"fb",x"f2",x"87"),
   114 => (x"38",x"33",x"32",x"4f"),
   115 => (x"53",x"44",x"41",x"44"),
   116 => (x"42",x"49",x"4e",x"00"),
   117 => (x"43",x"61",x"6e",x"27"),
   118 => (x"74",x"20",x"6c",x"6f"),
   119 => (x"61",x"64",x"20",x"66"),
   120 => (x"69",x"72",x"6d",x"77"),
   121 => (x"61",x"72",x"65",x"0a"),
   122 => (x"00",x"55",x"6e",x"61"),
   123 => (x"62",x"6c",x"65",x"20"),
   124 => (x"74",x"6f",x"20",x"6c"),
   125 => (x"6f",x"63",x"61",x"74"),
   126 => (x"65",x"20",x"70",x"61"),
   127 => (x"72",x"74",x"69",x"74"),
   128 => (x"69",x"6f",x"6e",x"0a"),
   129 => (x"00",x"48",x"75",x"6e"),
   130 => (x"74",x"69",x"6e",x"67"),
   131 => (x"20",x"66",x"6f",x"72"),
   132 => (x"20",x"70",x"61",x"72"),
   133 => (x"74",x"69",x"74",x"69"),
   134 => (x"6f",x"6e",x"0a",x"00"),
   135 => (x"49",x"6e",x"69",x"74"),
   136 => (x"69",x"61",x"6c",x"69"),
   137 => (x"7a",x"69",x"6e",x"67"),
   138 => (x"20",x"53",x"44",x"20"),
   139 => (x"63",x"61",x"72",x"64"),
   140 => (x"0a",x"00",x"46",x"61"),
   141 => (x"69",x"6c",x"65",x"64"),
   142 => (x"20",x"74",x"6f",x"20"),
   143 => (x"69",x"6e",x"69",x"74"),
   144 => (x"69",x"61",x"6c",x"69"),
   145 => (x"7a",x"65",x"20",x"53"),
   146 => (x"44",x"20",x"63",x"61"),
   147 => (x"72",x"64",x"0a",x"00"),
   148 => (x"00",x"00",x"00",x"00"),
   149 => (x"00",x"00",x"00",x"08"),
   150 => (x"33",x"fc",x"0f",x"ff"),
   151 => (x"00",x"df",x"f1",x"80"),
   152 => (x"60",x"f6",x"00",x"00"),
   153 => (x"00",x"12",x"1e",x"e4"),
   154 => (x"86",x"e3",x"48",x"c3"),
   155 => (x"ff",x"50",x"e3",x"97"),
   156 => (x"bf",x"7e",x"6e",x"49"),
   157 => (x"c3",x"ff",x"99",x"e3"),
   158 => (x"48",x"c3",x"ff",x"50"),
   159 => (x"c8",x"31",x"e3",x"97"),
   160 => (x"bf",x"48",x"c8",x"a6"),
   161 => (x"58",x"c3",x"ff",x"98"),
   162 => (x"cc",x"a6",x"58",x"70"),
   163 => (x"b1",x"e3",x"48",x"c3"),
   164 => (x"ff",x"50",x"c8",x"31"),
   165 => (x"e3",x"97",x"bf",x"48"),
   166 => (x"d0",x"a6",x"58",x"c3"),
   167 => (x"ff",x"98",x"d4",x"a6"),
   168 => (x"58",x"70",x"b1",x"e3"),
   169 => (x"48",x"c3",x"ff",x"50"),
   170 => (x"c8",x"31",x"e3",x"97"),
   171 => (x"bf",x"48",x"d8",x"a6"),
   172 => (x"58",x"c3",x"ff",x"98"),
   173 => (x"dc",x"a6",x"58",x"70"),
   174 => (x"b1",x"71",x"48",x"e4"),
   175 => (x"8e",x"26",x"4f",x"0e"),
   176 => (x"5e",x"5b",x"5c",x"0e"),
   177 => (x"1e",x"71",x"4a",x"49"),
   178 => (x"c3",x"ff",x"99",x"e3"),
   179 => (x"48",x"71",x"50",x"c1"),
   180 => (x"c0",x"ec",x"bf",x"05"),
   181 => (x"c8",x"87",x"d0",x"66"),
   182 => (x"48",x"c9",x"30",x"d4"),
   183 => (x"a6",x"58",x"d0",x"66"),
   184 => (x"49",x"d8",x"29",x"c3"),
   185 => (x"ff",x"99",x"e3",x"48"),
   186 => (x"71",x"50",x"d0",x"66"),
   187 => (x"49",x"d0",x"29",x"c3"),
   188 => (x"ff",x"99",x"e3",x"48"),
   189 => (x"71",x"50",x"d0",x"66"),
   190 => (x"49",x"c8",x"29",x"c3"),
   191 => (x"ff",x"99",x"e3",x"48"),
   192 => (x"71",x"50",x"d0",x"66"),
   193 => (x"49",x"c3",x"ff",x"99"),
   194 => (x"e3",x"48",x"71",x"50"),
   195 => (x"72",x"49",x"d0",x"29"),
   196 => (x"c3",x"ff",x"99",x"e3"),
   197 => (x"48",x"71",x"50",x"e3"),
   198 => (x"97",x"bf",x"7e",x"6e"),
   199 => (x"4b",x"c3",x"ff",x"9b"),
   200 => (x"c9",x"f0",x"ff",x"4c"),
   201 => (x"c3",x"ff",x"ab",x"05"),
   202 => (x"d9",x"87",x"e3",x"48"),
   203 => (x"c3",x"ff",x"50",x"e3"),
   204 => (x"97",x"bf",x"7e",x"6e"),
   205 => (x"4b",x"c3",x"ff",x"9b"),
   206 => (x"c1",x"8c",x"02",x"c6"),
   207 => (x"87",x"c3",x"ff",x"ab"),
   208 => (x"02",x"e7",x"87",x"73"),
   209 => (x"4a",x"c4",x"b7",x"2a"),
   210 => (x"c0",x"f0",x"a2",x"49"),
   211 => (x"c0",x"e6",x"cc",x"87"),
   212 => (x"73",x"4a",x"cf",x"9a"),
   213 => (x"c0",x"f0",x"a2",x"49"),
   214 => (x"c0",x"e6",x"c0",x"87"),
   215 => (x"73",x"48",x"26",x"c2"),
   216 => (x"87",x"26",x"4d",x"26"),
   217 => (x"4c",x"26",x"4b",x"26"),
   218 => (x"4f",x"1e",x"c0",x"49"),
   219 => (x"e3",x"48",x"c3",x"ff"),
   220 => (x"50",x"c1",x"81",x"c3"),
   221 => (x"c8",x"b7",x"a9",x"04"),
   222 => (x"f2",x"87",x"26",x"4f"),
   223 => (x"1e",x"73",x"1e",x"e8"),
   224 => (x"87",x"c4",x"f8",x"df"),
   225 => (x"4b",x"c0",x"1e",x"c0"),
   226 => (x"ff",x"f0",x"c1",x"f7"),
   227 => (x"49",x"fc",x"ef",x"87"),
   228 => (x"c4",x"86",x"c1",x"a8"),
   229 => (x"05",x"c0",x"e8",x"87"),
   230 => (x"e3",x"48",x"c3",x"ff"),
   231 => (x"50",x"c1",x"c0",x"c0"),
   232 => (x"c0",x"c0",x"c0",x"1e"),
   233 => (x"c0",x"e1",x"f0",x"c1"),
   234 => (x"e9",x"49",x"fc",x"d2"),
   235 => (x"87",x"c4",x"86",x"70"),
   236 => (x"98",x"05",x"c9",x"87"),
   237 => (x"e3",x"48",x"c3",x"ff"),
   238 => (x"50",x"c1",x"48",x"cb"),
   239 => (x"87",x"fe",x"e9",x"87"),
   240 => (x"c1",x"8b",x"05",x"fe"),
   241 => (x"ff",x"87",x"c0",x"48"),
   242 => (x"fe",x"da",x"87",x"1e"),
   243 => (x"73",x"1e",x"e3",x"48"),
   244 => (x"c3",x"ff",x"50",x"d0"),
   245 => (x"c5",x"49",x"c0",x"ef"),
   246 => (x"c7",x"87",x"d3",x"4b"),
   247 => (x"c0",x"1e",x"c0",x"ff"),
   248 => (x"f0",x"c1",x"c1",x"49"),
   249 => (x"fb",x"d8",x"87",x"c4"),
   250 => (x"86",x"70",x"98",x"05"),
   251 => (x"c9",x"87",x"e3",x"48"),
   252 => (x"c3",x"ff",x"50",x"c1"),
   253 => (x"48",x"cb",x"87",x"fd"),
   254 => (x"ef",x"87",x"c1",x"8b"),
   255 => (x"05",x"ff",x"dc",x"87"),
   256 => (x"c0",x"48",x"fd",x"e0"),
   257 => (x"87",x"43",x"6d",x"64"),
   258 => (x"5f",x"69",x"6e",x"69"),
   259 => (x"74",x"0a",x"00",x"1e"),
   260 => (x"73",x"1e",x"1e",x"fd"),
   261 => (x"d3",x"87",x"c6",x"ea"),
   262 => (x"1e",x"c0",x"e1",x"f0"),
   263 => (x"c1",x"c8",x"49",x"fa"),
   264 => (x"dd",x"87",x"70",x"4b"),
   265 => (x"1e",x"d2",x"fb",x"1e"),
   266 => (x"c0",x"ed",x"e1",x"87"),
   267 => (x"cc",x"86",x"c1",x"ab"),
   268 => (x"02",x"c8",x"87",x"fe"),
   269 => (x"d5",x"87",x"c0",x"48"),
   270 => (x"c1",x"fc",x"87",x"f8"),
   271 => (x"e8",x"87",x"70",x"49"),
   272 => (x"cf",x"ff",x"ff",x"99"),
   273 => (x"c6",x"ea",x"a9",x"02"),
   274 => (x"c8",x"87",x"fd",x"fe"),
   275 => (x"87",x"c0",x"48",x"c1"),
   276 => (x"e5",x"87",x"e3",x"48"),
   277 => (x"c3",x"ff",x"50",x"c0"),
   278 => (x"f1",x"4b",x"fc",x"df"),
   279 => (x"87",x"70",x"98",x"02"),
   280 => (x"c1",x"c3",x"87",x"c0"),
   281 => (x"1e",x"c0",x"ff",x"f0"),
   282 => (x"c1",x"fa",x"49",x"f9"),
   283 => (x"d1",x"87",x"c4",x"86"),
   284 => (x"70",x"98",x"05",x"c0"),
   285 => (x"f0",x"87",x"e3",x"48"),
   286 => (x"c3",x"ff",x"50",x"e3"),
   287 => (x"97",x"bf",x"7e",x"6e"),
   288 => (x"49",x"c3",x"ff",x"99"),
   289 => (x"e3",x"48",x"c3",x"ff"),
   290 => (x"50",x"e3",x"48",x"c3"),
   291 => (x"ff",x"50",x"e3",x"48"),
   292 => (x"c3",x"ff",x"50",x"e3"),
   293 => (x"48",x"c3",x"ff",x"50"),
   294 => (x"c1",x"c0",x"99",x"02"),
   295 => (x"c4",x"87",x"c1",x"48"),
   296 => (x"d5",x"87",x"c0",x"48"),
   297 => (x"d1",x"87",x"c2",x"ab"),
   298 => (x"05",x"c4",x"87",x"c0"),
   299 => (x"48",x"c8",x"87",x"c1"),
   300 => (x"8b",x"05",x"fe",x"e5"),
   301 => (x"87",x"c0",x"48",x"26"),
   302 => (x"fa",x"ea",x"87",x"63"),
   303 => (x"6d",x"64",x"5f",x"43"),
   304 => (x"4d",x"44",x"38",x"20"),
   305 => (x"72",x"65",x"73",x"70"),
   306 => (x"6f",x"6e",x"73",x"65"),
   307 => (x"3a",x"20",x"25",x"64"),
   308 => (x"0a",x"00",x"1e",x"73"),
   309 => (x"1e",x"c1",x"c0",x"ec"),
   310 => (x"48",x"c1",x"78",x"eb"),
   311 => (x"48",x"c3",x"ef",x"50"),
   312 => (x"c7",x"4b",x"e7",x"48"),
   313 => (x"c3",x"50",x"fa",x"c0"),
   314 => (x"87",x"e7",x"48",x"c2"),
   315 => (x"50",x"e3",x"48",x"c3"),
   316 => (x"ff",x"50",x"c0",x"1e"),
   317 => (x"c0",x"e5",x"d0",x"c1"),
   318 => (x"c0",x"49",x"f7",x"c2"),
   319 => (x"87",x"c4",x"86",x"c1"),
   320 => (x"a8",x"05",x"c1",x"87"),
   321 => (x"4b",x"c2",x"ab",x"05"),
   322 => (x"c5",x"87",x"c0",x"48"),
   323 => (x"c0",x"ef",x"87",x"c1"),
   324 => (x"8b",x"05",x"ff",x"cd"),
   325 => (x"87",x"fb",x"f7",x"87"),
   326 => (x"c1",x"c0",x"f0",x"58"),
   327 => (x"70",x"98",x"05",x"cd"),
   328 => (x"87",x"c1",x"1e",x"c0"),
   329 => (x"ff",x"f0",x"c1",x"d0"),
   330 => (x"49",x"f6",x"d3",x"87"),
   331 => (x"c4",x"86",x"e3",x"48"),
   332 => (x"c3",x"ff",x"50",x"e7"),
   333 => (x"48",x"c3",x"50",x"e3"),
   334 => (x"48",x"c3",x"ff",x"50"),
   335 => (x"c1",x"48",x"f8",x"e4"),
   336 => (x"87",x"0e",x"5e",x"5b"),
   337 => (x"5c",x"5d",x"0e",x"1e"),
   338 => (x"71",x"4a",x"c0",x"4d"),
   339 => (x"e3",x"48",x"c3",x"ff"),
   340 => (x"50",x"e7",x"48",x"c2"),
   341 => (x"50",x"eb",x"48",x"c7"),
   342 => (x"50",x"e3",x"48",x"c3"),
   343 => (x"ff",x"50",x"72",x"1e"),
   344 => (x"c0",x"ff",x"f0",x"c1"),
   345 => (x"d1",x"49",x"f5",x"d6"),
   346 => (x"87",x"c4",x"86",x"70"),
   347 => (x"98",x"05",x"c1",x"c5"),
   348 => (x"87",x"c5",x"ee",x"cd"),
   349 => (x"df",x"4b",x"e3",x"48"),
   350 => (x"c3",x"ff",x"50",x"e3"),
   351 => (x"97",x"bf",x"7e",x"6e"),
   352 => (x"49",x"c3",x"ff",x"99"),
   353 => (x"c3",x"fe",x"a9",x"05"),
   354 => (x"dd",x"87",x"c0",x"4c"),
   355 => (x"f3",x"d7",x"87",x"d4"),
   356 => (x"66",x"08",x"78",x"d4"),
   357 => (x"66",x"48",x"c4",x"80"),
   358 => (x"d8",x"a6",x"58",x"c1"),
   359 => (x"84",x"c2",x"c0",x"b7"),
   360 => (x"ac",x"04",x"e8",x"87"),
   361 => (x"c1",x"4b",x"4d",x"c1"),
   362 => (x"8b",x"05",x"ff",x"c9"),
   363 => (x"87",x"e3",x"48",x"c3"),
   364 => (x"ff",x"50",x"e7",x"48"),
   365 => (x"c3",x"50",x"75",x"48"),
   366 => (x"26",x"f6",x"e5",x"87"),
   367 => (x"1e",x"73",x"1e",x"71"),
   368 => (x"4b",x"49",x"d8",x"29"),
   369 => (x"c3",x"ff",x"99",x"73"),
   370 => (x"4a",x"c8",x"2a",x"cf"),
   371 => (x"fc",x"c0",x"9a",x"72"),
   372 => (x"b1",x"73",x"4a",x"c8"),
   373 => (x"32",x"c0",x"ff",x"f0"),
   374 => (x"c0",x"c0",x"9a",x"72"),
   375 => (x"b1",x"73",x"4a",x"d8"),
   376 => (x"32",x"ff",x"c0",x"c0"),
   377 => (x"c0",x"c0",x"9a",x"72"),
   378 => (x"b1",x"71",x"48",x"c4"),
   379 => (x"87",x"26",x"4d",x"26"),
   380 => (x"4c",x"26",x"4b",x"26"),
   381 => (x"4f",x"1e",x"73",x"1e"),
   382 => (x"71",x"4b",x"49",x"c8"),
   383 => (x"29",x"c3",x"ff",x"99"),
   384 => (x"73",x"4a",x"c8",x"32"),
   385 => (x"cf",x"fc",x"c0",x"9a"),
   386 => (x"72",x"b1",x"71",x"48"),
   387 => (x"e3",x"87",x"0e",x"5e"),
   388 => (x"5b",x"5c",x"0e",x"71"),
   389 => (x"4b",x"c0",x"4c",x"d0"),
   390 => (x"66",x"48",x"c0",x"b7"),
   391 => (x"a8",x"06",x"c0",x"e3"),
   392 => (x"87",x"13",x"4a",x"cc"),
   393 => (x"66",x"97",x"bf",x"49"),
   394 => (x"cc",x"66",x"48",x"c1"),
   395 => (x"80",x"d0",x"a6",x"58"),
   396 => (x"71",x"b7",x"aa",x"02"),
   397 => (x"c4",x"87",x"c1",x"48"),
   398 => (x"cc",x"87",x"c1",x"84"),
   399 => (x"d0",x"66",x"b7",x"ac"),
   400 => (x"04",x"ff",x"dd",x"87"),
   401 => (x"c0",x"48",x"c2",x"87"),
   402 => (x"26",x"4d",x"26",x"4c"),
   403 => (x"26",x"4b",x"26",x"4f"),
   404 => (x"0e",x"5e",x"5b",x"5c"),
   405 => (x"0e",x"1e",x"c1",x"c9"),
   406 => (x"e0",x"48",x"ff",x"78"),
   407 => (x"c1",x"c8",x"f8",x"48"),
   408 => (x"c0",x"78",x"c0",x"e6"),
   409 => (x"ec",x"49",x"c0",x"e4"),
   410 => (x"f7",x"87",x"c1",x"c0"),
   411 => (x"f0",x"1e",x"c0",x"49"),
   412 => (x"fb",x"ce",x"87",x"c4"),
   413 => (x"86",x"70",x"98",x"05"),
   414 => (x"c5",x"87",x"c0",x"48"),
   415 => (x"ca",x"e6",x"87",x"c0"),
   416 => (x"4b",x"c1",x"c9",x"dc"),
   417 => (x"48",x"c1",x"78",x"c8"),
   418 => (x"1e",x"c0",x"e6",x"f9"),
   419 => (x"1e",x"c1",x"c1",x"e6"),
   420 => (x"49",x"fd",x"fa",x"87"),
   421 => (x"c8",x"86",x"70",x"98"),
   422 => (x"05",x"c6",x"87",x"c1"),
   423 => (x"c9",x"dc",x"48",x"c0"),
   424 => (x"78",x"c8",x"1e",x"c0"),
   425 => (x"e7",x"c2",x"1e",x"c1"),
   426 => (x"c2",x"c2",x"49",x"fd"),
   427 => (x"e0",x"87",x"c8",x"86"),
   428 => (x"70",x"98",x"05",x"c6"),
   429 => (x"87",x"c1",x"c9",x"dc"),
   430 => (x"48",x"c0",x"78",x"c8"),
   431 => (x"1e",x"c0",x"e7",x"cb"),
   432 => (x"1e",x"c1",x"c2",x"c2"),
   433 => (x"49",x"fd",x"c6",x"87"),
   434 => (x"c8",x"86",x"70",x"98"),
   435 => (x"05",x"c5",x"87",x"c0"),
   436 => (x"48",x"c9",x"d1",x"87"),
   437 => (x"c1",x"c9",x"dc",x"bf"),
   438 => (x"1e",x"c0",x"e7",x"d4"),
   439 => (x"1e",x"c0",x"e2",x"ec"),
   440 => (x"87",x"c8",x"86",x"c1"),
   441 => (x"c9",x"dc",x"bf",x"02"),
   442 => (x"c1",x"ee",x"87",x"c1"),
   443 => (x"c0",x"f0",x"4a",x"48"),
   444 => (x"c6",x"fe",x"a0",x"4c"),
   445 => (x"c1",x"c7",x"f6",x"bf"),
   446 => (x"4b",x"c1",x"c8",x"ee"),
   447 => (x"9f",x"bf",x"49",x"72"),
   448 => (x"7e",x"c5",x"d6",x"ea"),
   449 => (x"a9",x"05",x"c0",x"cc"),
   450 => (x"87",x"c8",x"a4",x"4a"),
   451 => (x"6a",x"49",x"fa",x"eb"),
   452 => (x"87",x"70",x"4b",x"dc"),
   453 => (x"87",x"c7",x"fe",x"a2"),
   454 => (x"49",x"9f",x"69",x"49"),
   455 => (x"ca",x"e9",x"d5",x"a9"),
   456 => (x"02",x"c0",x"cd",x"87"),
   457 => (x"c0",x"e4",x"e9",x"49"),
   458 => (x"c0",x"e1",x"f5",x"87"),
   459 => (x"c0",x"48",x"c7",x"f4"),
   460 => (x"87",x"73",x"1e",x"c0"),
   461 => (x"e5",x"c7",x"1e",x"c0"),
   462 => (x"e1",x"d2",x"87",x"c1"),
   463 => (x"c0",x"f0",x"1e",x"73"),
   464 => (x"49",x"f7",x"fd",x"87"),
   465 => (x"cc",x"86",x"70",x"98"),
   466 => (x"05",x"c0",x"c5",x"87"),
   467 => (x"c0",x"48",x"c7",x"d4"),
   468 => (x"87",x"c0",x"e5",x"df"),
   469 => (x"49",x"c0",x"e1",x"c8"),
   470 => (x"87",x"c0",x"e7",x"e7"),
   471 => (x"1e",x"c0",x"e0",x"ec"),
   472 => (x"87",x"c8",x"1e",x"c0"),
   473 => (x"e7",x"ff",x"1e",x"c1"),
   474 => (x"c2",x"c2",x"49",x"fa"),
   475 => (x"e0",x"87",x"cc",x"86"),
   476 => (x"70",x"98",x"05",x"c0"),
   477 => (x"c9",x"87",x"c1",x"c8"),
   478 => (x"f8",x"48",x"c1",x"78"),
   479 => (x"c0",x"e3",x"87",x"c8"),
   480 => (x"1e",x"c0",x"e8",x"c8"),
   481 => (x"1e",x"c1",x"c1",x"e6"),
   482 => (x"49",x"fa",x"c2",x"87"),
   483 => (x"c8",x"86",x"70",x"98"),
   484 => (x"02",x"c0",x"ce",x"87"),
   485 => (x"c0",x"e6",x"c6",x"1e"),
   486 => (x"df",x"f2",x"87",x"c4"),
   487 => (x"86",x"c0",x"48",x"c6"),
   488 => (x"c3",x"87",x"c1",x"c8"),
   489 => (x"ee",x"97",x"bf",x"49"),
   490 => (x"c1",x"d5",x"a9",x"05"),
   491 => (x"c0",x"cd",x"87",x"c1"),
   492 => (x"c8",x"ef",x"97",x"bf"),
   493 => (x"49",x"c2",x"ea",x"a9"),
   494 => (x"02",x"c0",x"c5",x"87"),
   495 => (x"c0",x"48",x"c5",x"e4"),
   496 => (x"87",x"c1",x"c0",x"f0"),
   497 => (x"97",x"bf",x"49",x"c3"),
   498 => (x"e9",x"a9",x"02",x"c0"),
   499 => (x"d2",x"87",x"c1",x"c0"),
   500 => (x"f0",x"97",x"bf",x"49"),
   501 => (x"c3",x"eb",x"a9",x"02"),
   502 => (x"c0",x"c5",x"87",x"c0"),
   503 => (x"48",x"c5",x"c5",x"87"),
   504 => (x"c1",x"c0",x"fb",x"97"),
   505 => (x"bf",x"49",x"99",x"05"),
   506 => (x"c0",x"cc",x"87",x"c1"),
   507 => (x"c0",x"fc",x"97",x"bf"),
   508 => (x"49",x"c2",x"a9",x"02"),
   509 => (x"c0",x"c5",x"87",x"c0"),
   510 => (x"48",x"c4",x"e9",x"87"),
   511 => (x"c1",x"c0",x"fd",x"97"),
   512 => (x"bf",x"48",x"c1",x"c8"),
   513 => (x"f4",x"58",x"c1",x"88"),
   514 => (x"c1",x"c8",x"f8",x"58"),
   515 => (x"c1",x"c0",x"fe",x"97"),
   516 => (x"bf",x"49",x"73",x"81"),
   517 => (x"c1",x"c0",x"ff",x"97"),
   518 => (x"bf",x"4a",x"c8",x"32"),
   519 => (x"c1",x"c8",x"fc",x"48"),
   520 => (x"72",x"a1",x"78",x"c1"),
   521 => (x"c1",x"c0",x"97",x"bf"),
   522 => (x"48",x"c1",x"c9",x"d4"),
   523 => (x"58",x"c1",x"c8",x"f8"),
   524 => (x"bf",x"02",x"c2",x"e0"),
   525 => (x"87",x"c8",x"1e",x"c0"),
   526 => (x"e6",x"e3",x"1e",x"c1"),
   527 => (x"c2",x"c2",x"49",x"f7"),
   528 => (x"cc",x"87",x"c8",x"86"),
   529 => (x"70",x"98",x"02",x"c0"),
   530 => (x"c5",x"87",x"c0",x"48"),
   531 => (x"c3",x"d6",x"87",x"c1"),
   532 => (x"c8",x"f0",x"bf",x"48"),
   533 => (x"c4",x"30",x"c1",x"c9"),
   534 => (x"d8",x"58",x"c1",x"c8"),
   535 => (x"f0",x"bf",x"4a",x"c1"),
   536 => (x"c9",x"d0",x"5a",x"c1"),
   537 => (x"c1",x"d5",x"97",x"bf"),
   538 => (x"49",x"c8",x"31",x"c1"),
   539 => (x"c1",x"d4",x"97",x"bf"),
   540 => (x"4b",x"a1",x"49",x"c1"),
   541 => (x"c1",x"d6",x"97",x"bf"),
   542 => (x"4b",x"d0",x"33",x"73"),
   543 => (x"a1",x"49",x"c1",x"c1"),
   544 => (x"d7",x"97",x"bf",x"4b"),
   545 => (x"d8",x"33",x"73",x"a1"),
   546 => (x"49",x"c1",x"c9",x"dc"),
   547 => (x"59",x"c1",x"c9",x"d0"),
   548 => (x"bf",x"91",x"c1",x"c8"),
   549 => (x"fc",x"bf",x"81",x"c1"),
   550 => (x"c9",x"c4",x"59",x"c1"),
   551 => (x"c1",x"dd",x"97",x"bf"),
   552 => (x"4b",x"c8",x"33",x"c1"),
   553 => (x"c1",x"dc",x"97",x"bf"),
   554 => (x"4c",x"a3",x"4b",x"c1"),
   555 => (x"c1",x"de",x"97",x"bf"),
   556 => (x"4c",x"d0",x"34",x"74"),
   557 => (x"a3",x"4b",x"c1",x"c1"),
   558 => (x"df",x"97",x"bf",x"4c"),
   559 => (x"cf",x"9c",x"d8",x"34"),
   560 => (x"74",x"a3",x"4b",x"c1"),
   561 => (x"c9",x"c8",x"5b",x"c2"),
   562 => (x"8b",x"73",x"92",x"c1"),
   563 => (x"c9",x"c8",x"48",x"72"),
   564 => (x"a1",x"78",x"c1",x"ce"),
   565 => (x"87",x"c1",x"c1",x"c2"),
   566 => (x"97",x"bf",x"49",x"c8"),
   567 => (x"31",x"c1",x"c1",x"c1"),
   568 => (x"97",x"bf",x"4a",x"a1"),
   569 => (x"49",x"c1",x"c9",x"d8"),
   570 => (x"59",x"c5",x"31",x"c7"),
   571 => (x"ff",x"81",x"c9",x"29"),
   572 => (x"c1",x"c9",x"d0",x"59"),
   573 => (x"c1",x"c1",x"c7",x"97"),
   574 => (x"bf",x"4a",x"c8",x"32"),
   575 => (x"c1",x"c1",x"c6",x"97"),
   576 => (x"bf",x"4b",x"a2",x"4a"),
   577 => (x"c1",x"c9",x"dc",x"5a"),
   578 => (x"c1",x"c9",x"d0",x"bf"),
   579 => (x"92",x"c1",x"c8",x"fc"),
   580 => (x"bf",x"82",x"c1",x"c9"),
   581 => (x"cc",x"5a",x"c1",x"c9"),
   582 => (x"c4",x"48",x"c0",x"78"),
   583 => (x"c1",x"c9",x"c0",x"48"),
   584 => (x"72",x"a1",x"78",x"c1"),
   585 => (x"48",x"26",x"f4",x"e1"),
   586 => (x"87",x"4e",x"6f",x"20"),
   587 => (x"70",x"61",x"72",x"74"),
   588 => (x"69",x"74",x"69",x"6f"),
   589 => (x"6e",x"20",x"73",x"69"),
   590 => (x"67",x"6e",x"61",x"74"),
   591 => (x"75",x"72",x"65",x"20"),
   592 => (x"66",x"6f",x"75",x"6e"),
   593 => (x"64",x"0a",x"00",x"52"),
   594 => (x"65",x"61",x"64",x"69"),
   595 => (x"6e",x"67",x"20",x"62"),
   596 => (x"6f",x"6f",x"74",x"20"),
   597 => (x"73",x"65",x"63",x"74"),
   598 => (x"6f",x"72",x"20",x"25"),
   599 => (x"64",x"0a",x"00",x"52"),
   600 => (x"65",x"61",x"64",x"20"),
   601 => (x"62",x"6f",x"6f",x"74"),
   602 => (x"20",x"73",x"65",x"63"),
   603 => (x"74",x"6f",x"72",x"20"),
   604 => (x"66",x"72",x"6f",x"6d"),
   605 => (x"20",x"66",x"69",x"72"),
   606 => (x"73",x"74",x"20",x"70"),
   607 => (x"61",x"72",x"74",x"69"),
   608 => (x"74",x"69",x"6f",x"6e"),
   609 => (x"0a",x"00",x"55",x"6e"),
   610 => (x"73",x"75",x"70",x"70"),
   611 => (x"6f",x"72",x"74",x"65"),
   612 => (x"64",x"20",x"70",x"61"),
   613 => (x"72",x"74",x"69",x"74"),
   614 => (x"69",x"6f",x"6e",x"20"),
   615 => (x"74",x"79",x"70",x"65"),
   616 => (x"21",x"0d",x"00",x"46"),
   617 => (x"41",x"54",x"33",x"32"),
   618 => (x"20",x"20",x"20",x"00"),
   619 => (x"52",x"65",x"61",x"64"),
   620 => (x"69",x"6e",x"67",x"20"),
   621 => (x"4d",x"42",x"52",x"0a"),
   622 => (x"00",x"46",x"41",x"54"),
   623 => (x"31",x"36",x"20",x"20"),
   624 => (x"20",x"00",x"46",x"41"),
   625 => (x"54",x"33",x"32",x"20"),
   626 => (x"20",x"20",x"00",x"46"),
   627 => (x"41",x"54",x"31",x"32"),
   628 => (x"20",x"20",x"20",x"00"),
   629 => (x"50",x"61",x"72",x"74"),
   630 => (x"69",x"74",x"69",x"6f"),
   631 => (x"6e",x"63",x"6f",x"75"),
   632 => (x"6e",x"74",x"20",x"25"),
   633 => (x"64",x"0a",x"00",x"48"),
   634 => (x"75",x"6e",x"74",x"69"),
   635 => (x"6e",x"67",x"20",x"66"),
   636 => (x"6f",x"72",x"20",x"66"),
   637 => (x"69",x"6c",x"65",x"73"),
   638 => (x"79",x"73",x"74",x"65"),
   639 => (x"6d",x"0a",x"00",x"46"),
   640 => (x"41",x"54",x"33",x"32"),
   641 => (x"20",x"20",x"20",x"00"),
   642 => (x"46",x"41",x"54",x"31"),
   643 => (x"36",x"20",x"20",x"20"),
   644 => (x"00",x"0e",x"5e",x"5b"),
   645 => (x"5c",x"5d",x"0e",x"71"),
   646 => (x"4a",x"c1",x"c8",x"f8"),
   647 => (x"bf",x"02",x"cc",x"87"),
   648 => (x"72",x"4b",x"c7",x"b7"),
   649 => (x"2b",x"72",x"4c",x"c1"),
   650 => (x"ff",x"9c",x"ca",x"87"),
   651 => (x"72",x"4b",x"c8",x"b7"),
   652 => (x"2b",x"72",x"4c",x"c3"),
   653 => (x"ff",x"9c",x"c1",x"c9"),
   654 => (x"e0",x"bf",x"ab",x"02"),
   655 => (x"de",x"87",x"c1",x"c0"),
   656 => (x"f0",x"1e",x"c1",x"c8"),
   657 => (x"fc",x"bf",x"49",x"73"),
   658 => (x"81",x"eb",x"f5",x"87"),
   659 => (x"c4",x"86",x"70",x"98"),
   660 => (x"05",x"c5",x"87",x"c0"),
   661 => (x"48",x"c0",x"f5",x"87"),
   662 => (x"c1",x"c9",x"e4",x"5b"),
   663 => (x"c1",x"c8",x"f8",x"bf"),
   664 => (x"02",x"d8",x"87",x"74"),
   665 => (x"4a",x"c4",x"92",x"c1"),
   666 => (x"c0",x"f0",x"82",x"6a"),
   667 => (x"49",x"ed",x"cc",x"87"),
   668 => (x"70",x"49",x"4d",x"cf"),
   669 => (x"ff",x"ff",x"ff",x"ff"),
   670 => (x"9d",x"d0",x"87",x"74"),
   671 => (x"4a",x"c2",x"92",x"c1"),
   672 => (x"c0",x"f0",x"82",x"9f"),
   673 => (x"6a",x"49",x"ed",x"ec"),
   674 => (x"87",x"70",x"4d",x"75"),
   675 => (x"48",x"ee",x"f8",x"87"),
   676 => (x"0e",x"5e",x"5b",x"5c"),
   677 => (x"5d",x"0e",x"f4",x"86"),
   678 => (x"71",x"4c",x"c0",x"4b"),
   679 => (x"c1",x"c9",x"e0",x"48"),
   680 => (x"ff",x"78",x"c1",x"c9"),
   681 => (x"c4",x"bf",x"4d",x"c1"),
   682 => (x"c9",x"c8",x"bf",x"7e"),
   683 => (x"c1",x"c8",x"f8",x"bf"),
   684 => (x"02",x"c9",x"87",x"c1"),
   685 => (x"c8",x"f0",x"bf",x"4a"),
   686 => (x"c4",x"32",x"c7",x"87"),
   687 => (x"c1",x"c9",x"cc",x"bf"),
   688 => (x"4a",x"c4",x"32",x"c8"),
   689 => (x"a6",x"5a",x"c8",x"a6"),
   690 => (x"48",x"c0",x"78",x"c4"),
   691 => (x"66",x"48",x"c0",x"a8"),
   692 => (x"06",x"c3",x"cc",x"87"),
   693 => (x"c8",x"66",x"49",x"cf"),
   694 => (x"99",x"05",x"c0",x"e2"),
   695 => (x"87",x"6e",x"1e",x"c0"),
   696 => (x"ef",x"e1",x"1e",x"d2"),
   697 => (x"e7",x"87",x"c1",x"c0"),
   698 => (x"f0",x"1e",x"cc",x"66"),
   699 => (x"49",x"48",x"c1",x"80"),
   700 => (x"d0",x"a6",x"58",x"71"),
   701 => (x"e9",x"ca",x"87",x"cc"),
   702 => (x"86",x"c1",x"c0",x"f0"),
   703 => (x"4b",x"c3",x"87",x"c0"),
   704 => (x"e0",x"83",x"97",x"6b"),
   705 => (x"49",x"99",x"02",x"c2"),
   706 => (x"c4",x"87",x"97",x"6b"),
   707 => (x"49",x"c3",x"e5",x"a9"),
   708 => (x"02",x"c1",x"fa",x"87"),
   709 => (x"cb",x"a3",x"49",x"97"),
   710 => (x"69",x"49",x"d8",x"99"),
   711 => (x"05",x"c1",x"ee",x"87"),
   712 => (x"cb",x"1e",x"c0",x"e0"),
   713 => (x"66",x"1e",x"73",x"49"),
   714 => (x"eb",x"e3",x"87",x"c8"),
   715 => (x"86",x"70",x"98",x"05"),
   716 => (x"c1",x"db",x"87",x"dc"),
   717 => (x"a3",x"4a",x"6a",x"49"),
   718 => (x"ea",x"c1",x"87",x"70"),
   719 => (x"4a",x"c4",x"a4",x"49"),
   720 => (x"72",x"79",x"da",x"a3"),
   721 => (x"4a",x"9f",x"6a",x"49"),
   722 => (x"ea",x"ea",x"87",x"70"),
   723 => (x"7e",x"c1",x"c8",x"f8"),
   724 => (x"bf",x"02",x"d8",x"87"),
   725 => (x"d4",x"a3",x"4a",x"9f"),
   726 => (x"6a",x"49",x"ea",x"d8"),
   727 => (x"87",x"70",x"49",x"c0"),
   728 => (x"ff",x"ff",x"99",x"71"),
   729 => (x"48",x"d0",x"30",x"c8"),
   730 => (x"a6",x"58",x"c5",x"87"),
   731 => (x"c4",x"a6",x"48",x"c0"),
   732 => (x"78",x"c4",x"66",x"4a"),
   733 => (x"6e",x"82",x"c8",x"a4"),
   734 => (x"49",x"72",x"79",x"c0"),
   735 => (x"7c",x"dc",x"66",x"1e"),
   736 => (x"c0",x"ef",x"fe",x"1e"),
   737 => (x"d0",x"c6",x"87",x"c8"),
   738 => (x"86",x"c1",x"48",x"c1"),
   739 => (x"ce",x"87",x"c8",x"66"),
   740 => (x"48",x"c1",x"80",x"cc"),
   741 => (x"a6",x"58",x"c8",x"66"),
   742 => (x"48",x"c4",x"66",x"a8"),
   743 => (x"04",x"fc",x"f4",x"87"),
   744 => (x"c1",x"c8",x"f8",x"bf"),
   745 => (x"02",x"c0",x"f2",x"87"),
   746 => (x"75",x"49",x"f9",x"e4"),
   747 => (x"87",x"70",x"4d",x"1e"),
   748 => (x"c0",x"f0",x"cf",x"1e"),
   749 => (x"cf",x"d6",x"87",x"c8"),
   750 => (x"86",x"75",x"49",x"cf"),
   751 => (x"ff",x"ff",x"ff",x"f8"),
   752 => (x"99",x"a9",x"02",x"d5"),
   753 => (x"87",x"75",x"49",x"c2"),
   754 => (x"89",x"c1",x"c8",x"f0"),
   755 => (x"bf",x"91",x"c1",x"c9"),
   756 => (x"c0",x"bf",x"48",x"71"),
   757 => (x"80",x"70",x"7e",x"fb"),
   758 => (x"ec",x"87",x"c0",x"48"),
   759 => (x"f4",x"8e",x"e9",x"e7"),
   760 => (x"87",x"52",x"65",x"61"),
   761 => (x"64",x"69",x"6e",x"67"),
   762 => (x"20",x"64",x"69",x"72"),
   763 => (x"65",x"63",x"74",x"6f"),
   764 => (x"72",x"79",x"20",x"73"),
   765 => (x"65",x"63",x"74",x"6f"),
   766 => (x"72",x"20",x"25",x"64"),
   767 => (x"0a",x"00",x"66",x"69"),
   768 => (x"6c",x"65",x"20",x"22"),
   769 => (x"25",x"73",x"22",x"20"),
   770 => (x"66",x"6f",x"75",x"6e"),
   771 => (x"64",x"0d",x"00",x"47"),
   772 => (x"65",x"74",x"46",x"41"),
   773 => (x"54",x"4c",x"69",x"6e"),
   774 => (x"6b",x"20",x"72",x"65"),
   775 => (x"74",x"75",x"72",x"6e"),
   776 => (x"65",x"64",x"20",x"25"),
   777 => (x"64",x"0a",x"00",x"0e"),
   778 => (x"5e",x"5b",x"5c",x"5d"),
   779 => (x"0e",x"1e",x"71",x"4b"),
   780 => (x"1e",x"c1",x"c9",x"e4"),
   781 => (x"49",x"f9",x"d8",x"87"),
   782 => (x"c4",x"86",x"70",x"98"),
   783 => (x"02",x"c1",x"f5",x"87"),
   784 => (x"c1",x"c9",x"e8",x"bf"),
   785 => (x"49",x"c7",x"ff",x"81"),
   786 => (x"c9",x"29",x"71",x"7e"),
   787 => (x"c0",x"4d",x"4c",x"6e"),
   788 => (x"48",x"c0",x"b7",x"a8"),
   789 => (x"06",x"c1",x"ec",x"87"),
   790 => (x"c1",x"c9",x"c0",x"bf"),
   791 => (x"49",x"c1",x"c9",x"ec"),
   792 => (x"bf",x"4a",x"c2",x"8a"),
   793 => (x"c1",x"c8",x"f0",x"bf"),
   794 => (x"92",x"72",x"a1",x"49"),
   795 => (x"c1",x"c8",x"f4",x"bf"),
   796 => (x"4a",x"74",x"9a",x"72"),
   797 => (x"a1",x"49",x"d4",x"66"),
   798 => (x"1e",x"71",x"e3",x"c4"),
   799 => (x"87",x"c4",x"86",x"70"),
   800 => (x"98",x"05",x"c5",x"87"),
   801 => (x"c0",x"48",x"c1",x"c0"),
   802 => (x"87",x"c1",x"84",x"c1"),
   803 => (x"c8",x"f4",x"bf",x"49"),
   804 => (x"74",x"99",x"05",x"cc"),
   805 => (x"87",x"c1",x"c9",x"ec"),
   806 => (x"bf",x"49",x"f5",x"f4"),
   807 => (x"87",x"c1",x"c9",x"f0"),
   808 => (x"58",x"d4",x"66",x"48"),
   809 => (x"c8",x"c0",x"80",x"d8"),
   810 => (x"a6",x"58",x"c1",x"85"),
   811 => (x"6e",x"b7",x"ad",x"04"),
   812 => (x"fe",x"e5",x"87",x"cf"),
   813 => (x"87",x"73",x"1e",x"c0"),
   814 => (x"f3",x"cd",x"1e",x"cb"),
   815 => (x"cf",x"87",x"c8",x"86"),
   816 => (x"c0",x"48",x"c5",x"87"),
   817 => (x"c1",x"c9",x"e8",x"bf"),
   818 => (x"48",x"26",x"e5",x"fb"),
   819 => (x"87",x"43",x"61",x"6e"),
   820 => (x"27",x"74",x"20",x"6f"),
   821 => (x"70",x"65",x"6e",x"20"),
   822 => (x"25",x"73",x"0a",x"00"),
   823 => (x"1e",x"f3",x"48",x"71"),
   824 => (x"50",x"48",x"26",x"4f"),
   825 => (x"0e",x"5e",x"5b",x"5c"),
   826 => (x"5d",x"0e",x"f8",x"86"),
   827 => (x"71",x"4a",x"c0",x"e4"),
   828 => (x"66",x"4c",x"d5",x"fb"),
   829 => (x"a7",x"4b",x"c2",x"cb"),
   830 => (x"a7",x"7e",x"c4",x"a6"),
   831 => (x"48",x"c0",x"78",x"72"),
   832 => (x"9a",x"05",x"c6",x"87"),
   833 => (x"c0",x"f0",x"53",x"c1"),
   834 => (x"c7",x"87",x"72",x"9a"),
   835 => (x"02",x"c0",x"e3",x"87"),
   836 => (x"d8",x"66",x"4d",x"72"),
   837 => (x"1e",x"72",x"49",x"75"),
   838 => (x"4a",x"ca",x"e9",x"87"),
   839 => (x"26",x"4a",x"6e",x"81"),
   840 => (x"11",x"53",x"72",x"49"),
   841 => (x"75",x"4a",x"ca",x"dc"),
   842 => (x"87",x"70",x"4a",x"c1"),
   843 => (x"8c",x"72",x"9a",x"05"),
   844 => (x"ff",x"e0",x"87",x"c0"),
   845 => (x"b7",x"ac",x"06",x"d8"),
   846 => (x"87",x"c0",x"e8",x"66"),
   847 => (x"02",x"c5",x"87",x"c0"),
   848 => (x"f0",x"4a",x"c3",x"87"),
   849 => (x"c0",x"e0",x"4a",x"72"),
   850 => (x"53",x"c1",x"8c",x"c0"),
   851 => (x"b7",x"ac",x"01",x"e8"),
   852 => (x"87",x"d4",x"dc",x"a7"),
   853 => (x"ab",x"02",x"df",x"87"),
   854 => (x"dc",x"66",x"4c",x"c0"),
   855 => (x"e0",x"66",x"1e",x"c1"),
   856 => (x"8b",x"97",x"6b",x"49"),
   857 => (x"74",x"0f",x"c4",x"86"),
   858 => (x"66",x"48",x"c1",x"80"),
   859 => (x"c8",x"a6",x"58",x"d3"),
   860 => (x"fe",x"a7",x"ab",x"05"),
   861 => (x"ff",x"e4",x"87",x"c4"),
   862 => (x"66",x"48",x"f8",x"8e"),
   863 => (x"26",x"4d",x"26",x"4c"),
   864 => (x"26",x"4b",x"26",x"4f"),
   865 => (x"30",x"31",x"32",x"33"),
   866 => (x"34",x"35",x"36",x"37"),
   867 => (x"38",x"39",x"41",x"42"),
   868 => (x"43",x"44",x"45",x"46"),
   869 => (x"00",x"0e",x"5e",x"5b"),
   870 => (x"5c",x"5d",x"0e",x"71"),
   871 => (x"4b",x"ff",x"4d",x"13"),
   872 => (x"4c",x"9c",x"02",x"d7"),
   873 => (x"87",x"c1",x"85",x"d4"),
   874 => (x"66",x"1e",x"74",x"49"),
   875 => (x"d4",x"66",x"0f",x"c4"),
   876 => (x"86",x"74",x"a8",x"05"),
   877 => (x"c6",x"87",x"13",x"4c"),
   878 => (x"9c",x"05",x"e9",x"87"),
   879 => (x"75",x"48",x"26",x"4d"),
   880 => (x"26",x"4c",x"26",x"4b"),
   881 => (x"26",x"4f",x"0e",x"5e"),
   882 => (x"5b",x"5c",x"5d",x"0e"),
   883 => (x"e8",x"86",x"c8",x"a6"),
   884 => (x"59",x"c0",x"e8",x"66"),
   885 => (x"4d",x"c0",x"4c",x"c8"),
   886 => (x"a6",x"48",x"c0",x"78"),
   887 => (x"c4",x"66",x"97",x"bf"),
   888 => (x"4b",x"c4",x"66",x"48"),
   889 => (x"c1",x"80",x"c8",x"a6"),
   890 => (x"58",x"73",x"9b",x"02"),
   891 => (x"c6",x"d2",x"87",x"c8"),
   892 => (x"66",x"02",x"c5",x"d8"),
   893 => (x"87",x"cc",x"a6",x"48"),
   894 => (x"c0",x"78",x"fc",x"80"),
   895 => (x"c0",x"78",x"73",x"4a"),
   896 => (x"c0",x"e0",x"8a",x"02"),
   897 => (x"c3",x"c8",x"87",x"c3"),
   898 => (x"8a",x"02",x"c3",x"c2"),
   899 => (x"87",x"c2",x"8a",x"02"),
   900 => (x"c2",x"ea",x"87",x"8a"),
   901 => (x"02",x"c2",x"f7",x"87"),
   902 => (x"c4",x"8a",x"02",x"c2"),
   903 => (x"f1",x"87",x"c2",x"8a"),
   904 => (x"02",x"c2",x"eb",x"87"),
   905 => (x"c3",x"8a",x"02",x"c2"),
   906 => (x"ed",x"87",x"d4",x"8a"),
   907 => (x"02",x"c0",x"fa",x"87"),
   908 => (x"8a",x"02",x"c1",x"c5"),
   909 => (x"87",x"ca",x"8a",x"02"),
   910 => (x"c0",x"f7",x"87",x"c1"),
   911 => (x"8a",x"02",x"c1",x"e5"),
   912 => (x"87",x"8a",x"02",x"c0"),
   913 => (x"e4",x"87",x"c5",x"8a"),
   914 => (x"02",x"df",x"87",x"c3"),
   915 => (x"8a",x"02",x"c1",x"cd"),
   916 => (x"87",x"c4",x"8a",x"02"),
   917 => (x"c0",x"e3",x"87",x"c3"),
   918 => (x"8a",x"02",x"c0",x"e5"),
   919 => (x"87",x"c2",x"8a",x"02"),
   920 => (x"c8",x"87",x"c3",x"8a"),
   921 => (x"02",x"d3",x"87",x"c1"),
   922 => (x"f9",x"87",x"cc",x"a6"),
   923 => (x"48",x"ca",x"78",x"c2"),
   924 => (x"d2",x"87",x"cc",x"a6"),
   925 => (x"48",x"c2",x"78",x"c2"),
   926 => (x"ca",x"87",x"cc",x"a6"),
   927 => (x"48",x"d0",x"78",x"c2"),
   928 => (x"c2",x"87",x"c0",x"f0"),
   929 => (x"66",x"1e",x"c0",x"f0"),
   930 => (x"66",x"1e",x"c4",x"85"),
   931 => (x"75",x"4a",x"c4",x"8a"),
   932 => (x"6a",x"49",x"fc",x"c0"),
   933 => (x"87",x"c8",x"86",x"70"),
   934 => (x"49",x"a4",x"4c",x"c1"),
   935 => (x"e6",x"87",x"c8",x"a6"),
   936 => (x"48",x"c1",x"78",x"c1"),
   937 => (x"de",x"87",x"c0",x"f0"),
   938 => (x"66",x"1e",x"c4",x"85"),
   939 => (x"75",x"4a",x"c4",x"8a"),
   940 => (x"6a",x"49",x"c0",x"f0"),
   941 => (x"66",x"0f",x"c4",x"86"),
   942 => (x"c1",x"84",x"c1",x"c7"),
   943 => (x"87",x"c0",x"f0",x"66"),
   944 => (x"1e",x"c0",x"e5",x"49"),
   945 => (x"c0",x"f0",x"66",x"0f"),
   946 => (x"c4",x"86",x"c1",x"84"),
   947 => (x"c0",x"f5",x"87",x"c8"),
   948 => (x"a6",x"48",x"c1",x"78"),
   949 => (x"c0",x"ed",x"87",x"d0"),
   950 => (x"a6",x"48",x"c1",x"78"),
   951 => (x"f8",x"80",x"c1",x"78"),
   952 => (x"c0",x"e1",x"87",x"c0"),
   953 => (x"f0",x"ab",x"06",x"db"),
   954 => (x"87",x"c0",x"f9",x"ab"),
   955 => (x"03",x"d5",x"87",x"d4"),
   956 => (x"66",x"49",x"ca",x"91"),
   957 => (x"73",x"4a",x"c0",x"f0"),
   958 => (x"8a",x"d4",x"a6",x"48"),
   959 => (x"72",x"a1",x"78",x"c8"),
   960 => (x"a6",x"48",x"c1",x"78"),
   961 => (x"cc",x"66",x"02",x"c1"),
   962 => (x"e4",x"87",x"c4",x"85"),
   963 => (x"75",x"49",x"c4",x"89"),
   964 => (x"69",x"7e",x"c1",x"e4"),
   965 => (x"ab",x"05",x"d5",x"87"),
   966 => (x"6e",x"48",x"c0",x"b7"),
   967 => (x"a8",x"03",x"cd",x"87"),
   968 => (x"c0",x"ed",x"49",x"f6"),
   969 => (x"f6",x"87",x"6e",x"48"),
   970 => (x"c0",x"08",x"88",x"70"),
   971 => (x"7e",x"d0",x"66",x"1e"),
   972 => (x"d8",x"66",x"1e",x"c0"),
   973 => (x"f8",x"66",x"1e",x"c0"),
   974 => (x"f8",x"66",x"1e",x"dc"),
   975 => (x"66",x"1e",x"d4",x"66"),
   976 => (x"49",x"f6",x"e0",x"87"),
   977 => (x"d4",x"86",x"70",x"49"),
   978 => (x"a4",x"4c",x"c0",x"e1"),
   979 => (x"87",x"c0",x"e5",x"ab"),
   980 => (x"05",x"cf",x"87",x"d0"),
   981 => (x"a6",x"48",x"c0",x"78"),
   982 => (x"c4",x"80",x"c0",x"78"),
   983 => (x"f4",x"80",x"c1",x"78"),
   984 => (x"cc",x"87",x"c0",x"f0"),
   985 => (x"66",x"1e",x"73",x"49"),
   986 => (x"c0",x"f0",x"66",x"0f"),
   987 => (x"c4",x"86",x"c4",x"66"),
   988 => (x"97",x"bf",x"4b",x"c4"),
   989 => (x"66",x"48",x"c1",x"80"),
   990 => (x"c8",x"a6",x"58",x"73"),
   991 => (x"9b",x"05",x"f9",x"ee"),
   992 => (x"87",x"74",x"48",x"e8"),
   993 => (x"8e",x"26",x"4d",x"26"),
   994 => (x"4c",x"26",x"4b",x"26"),
   995 => (x"4f",x"1e",x"c0",x"1e"),
   996 => (x"f5",x"c9",x"a7",x"1e"),
   997 => (x"d0",x"a6",x"1e",x"d0"),
   998 => (x"66",x"49",x"f8",x"e9"),
   999 => (x"87",x"f4",x"8e",x"26"),
  1000 => (x"4f",x"0e",x"5e",x"5b"),
  1001 => (x"5c",x"0e",x"71",x"4b"),
  1002 => (x"c0",x"4c",x"13",x"4a"),
  1003 => (x"9a",x"02",x"cd",x"87"),
  1004 => (x"72",x"49",x"f4",x"e7"),
  1005 => (x"87",x"c1",x"84",x"13"),
  1006 => (x"4a",x"9a",x"05",x"f3"),
  1007 => (x"87",x"74",x"48",x"26"),
  1008 => (x"4c",x"26",x"4b",x"26"),
  1009 => (x"4f",x"1e",x"73",x"1e"),
  1010 => (x"72",x"9a",x"02",x"c0"),
  1011 => (x"e7",x"87",x"c0",x"48"),
  1012 => (x"c1",x"4b",x"72",x"a9"),
  1013 => (x"06",x"d1",x"87",x"72"),
  1014 => (x"82",x"06",x"c9",x"87"),
  1015 => (x"73",x"83",x"72",x"a9"),
  1016 => (x"01",x"f4",x"87",x"c3"),
  1017 => (x"87",x"c1",x"b2",x"3a"),
  1018 => (x"72",x"a9",x"03",x"89"),
  1019 => (x"73",x"80",x"07",x"c1"),
  1020 => (x"2a",x"2b",x"05",x"f3"),
  1021 => (x"87",x"26",x"4b",x"26"),
  1022 => (x"4f",x"1e",x"75",x"1e"),
  1023 => (x"c4",x"4d",x"71",x"b7"),
  1024 => (x"a1",x"04",x"ff",x"b9"),
  1025 => (x"c1",x"81",x"c3",x"bd"),
  1026 => (x"07",x"72",x"b7",x"a2"),
  1027 => (x"04",x"ff",x"ba",x"c1"),
  1028 => (x"82",x"c1",x"bd",x"07"),
  1029 => (x"fe",x"ee",x"87",x"c1"),
  1030 => (x"2d",x"04",x"ff",x"b8"),
  1031 => (x"c1",x"80",x"07",x"2d"),
  1032 => (x"04",x"ff",x"b9",x"c1"),
  1033 => (x"81",x"07",x"26",x"4d"),
  1034 => (x"26",x"4f",x"26",x"4d"),
	others => (others => x"00")
);

-- Xilinx XST attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "no_rw_check";

-- Altera Quartus attributes
attribute ramstyle: string;
attribute ramstyle of ram: signal is "no_rw_check";

signal q_local : word_t;
signal q2_local : word_t;

begin
    
	process(clk,q_local)
	begin

		q(31 downto 24)<=q_local(0);
		q(23 downto 16)<=q_local(1);
		q(15 downto 8)<=q_local(2);
		q(7 downto 0)<=q_local(3);

		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel(3) = '1') then
					ram(to_integer(unsigned(addr)))(3) <= d(7 downto 0);
				end if;
				if bytesel(2) = '1' then
					ram(to_integer(unsigned(addr)))(2) <= d(15 downto 8);
				end if;
				if bytesel(1) = '1' then
					ram(to_integer(unsigned(addr)))(1) <= d(23 downto 16);
				end if;
				if bytesel(0) = '1' then
					ram(to_integer(unsigned(addr)))(0) <= d(31 downto 24);
				end if;
			end if;
			q_local <= ram(to_integer(unsigned(addr)));
		end if;
	end process;

	-- Second port
	
	process(clk,q2_local)
	begin

		q2(31 downto 24)<=q2_local(0);
		q2(23 downto 16)<=q2_local(1);
		q2(15 downto 8)<=q2_local(2);
		q2(7 downto 0)<=q2_local(3);

		if(rising_edge(clk)) then 
			if(we2 = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel2(3) = '1') then
					ram(to_integer(unsigned(addr2)))(3) <= d2(7 downto 0);
				end if;
				if bytesel2(2) = '1' then
					ram(to_integer(unsigned(addr2)))(2) <= d2(15 downto 8);
				end if;
				if bytesel2(1) = '1' then
					ram(to_integer(unsigned(addr2)))(1) <= d2(23 downto 16);
				end if;
				if bytesel2(0) = '1' then
					ram(to_integer(unsigned(addr2)))(0) <= d2(31 downto 24);
				end if;
			end if;
			q2_local <= ram(to_integer(unsigned(addr2)));
		end if;
	end process;

end arch;

