library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"01",
     1 => x"da",
     2 => x"87",
     3 => x"04",
     4 => x"dd",
     5 => x"87",
     6 => x"0e",
     7 => x"58",
     8 => x"5e",
     9 => x"59",
    10 => x"5a",
    11 => x"0e",
    12 => x"27",
    13 => x"00",
    14 => x"00",
    15 => x"00",
    16 => x"2c",
    17 => x"0f",
    18 => x"26",
    19 => x"4a",
    20 => x"26",
    21 => x"49",
    22 => x"26",
    23 => x"48",
    24 => x"ff",
    25 => x"80",
    26 => x"26",
    27 => x"08",
    28 => x"4f",
    29 => x"27",
    30 => x"00",
    31 => x"00",
    32 => x"00",
    33 => x"2d",
    34 => x"4f",
    35 => x"27",
    36 => x"00",
    37 => x"00",
    38 => x"00",
    39 => x"29",
    40 => x"4f",
    41 => x"00",
    42 => x"fd",
    43 => x"87",
    44 => x"4f",
    45 => x"c1",
    46 => x"d1",
    47 => x"ec",
    48 => x"4e",
    49 => x"c9",
    50 => x"c0",
    51 => x"86",
    52 => x"c1",
    53 => x"d1",
    54 => x"ec",
    55 => x"49",
    56 => x"c1",
    57 => x"c7",
    58 => x"e8",
    59 => x"48",
    60 => x"89",
    61 => x"d0",
    62 => x"89",
    63 => x"03",
    64 => x"c0",
    65 => x"40",
    66 => x"40",
    67 => x"40",
    68 => x"40",
    69 => x"f6",
    70 => x"87",
    71 => x"d0",
    72 => x"81",
    73 => x"05",
    74 => x"c0",
    75 => x"50",
    76 => x"c1",
    77 => x"89",
    78 => x"05",
    79 => x"f9",
    80 => x"87",
    81 => x"c1",
    82 => x"c7",
    83 => x"e8",
    84 => x"4d",
    85 => x"c1",
    86 => x"c7",
    87 => x"e8",
    88 => x"4c",
    89 => x"74",
    90 => x"ad",
    91 => x"02",
    92 => x"c4",
    93 => x"87",
    94 => x"24",
    95 => x"0f",
    96 => x"f7",
    97 => x"87",
    98 => x"c1",
    99 => x"e3",
   100 => x"87",
   101 => x"c1",
   102 => x"c7",
   103 => x"e8",
   104 => x"4d",
   105 => x"c1",
   106 => x"c7",
   107 => x"e8",
   108 => x"4c",
   109 => x"74",
   110 => x"ad",
   111 => x"02",
   112 => x"c6",
   113 => x"87",
   114 => x"c4",
   115 => x"8c",
   116 => x"6c",
   117 => x"0f",
   118 => x"f5",
   119 => x"87",
   120 => x"00",
   121 => x"fd",
   122 => x"87",
   123 => x"1e",
   124 => x"73",
   125 => x"1e",
   126 => x"c2",
   127 => x"c0",
   128 => x"c0",
   129 => x"4b",
   130 => x"73",
   131 => x"0f",
   132 => x"c4",
   133 => x"87",
   134 => x"26",
   135 => x"4d",
   136 => x"26",
   137 => x"4c",
   138 => x"26",
   139 => x"4b",
   140 => x"26",
   141 => x"4f",
   142 => x"0e",
   143 => x"5e",
   144 => x"5b",
   145 => x"5c",
   146 => x"0e",
   147 => x"71",
   148 => x"4a",
   149 => x"c0",
   150 => x"4c",
   151 => x"72",
   152 => x"4b",
   153 => x"dc",
   154 => x"b7",
   155 => x"2b",
   156 => x"cf",
   157 => x"9b",
   158 => x"c4",
   159 => x"32",
   160 => x"c9",
   161 => x"b7",
   162 => x"ab",
   163 => x"06",
   164 => x"c5",
   165 => x"87",
   166 => x"c0",
   167 => x"f7",
   168 => x"83",
   169 => x"c3",
   170 => x"87",
   171 => x"c0",
   172 => x"f0",
   173 => x"83",
   174 => x"cc",
   175 => x"66",
   176 => x"0b",
   177 => x"97",
   178 => x"7b",
   179 => x"0b",
   180 => x"cc",
   181 => x"66",
   182 => x"48",
   183 => x"c1",
   184 => x"80",
   185 => x"d0",
   186 => x"a6",
   187 => x"58",
   188 => x"c1",
   189 => x"84",
   190 => x"c8",
   191 => x"b7",
   192 => x"ac",
   193 => x"04",
   194 => x"ff",
   195 => x"d2",
   196 => x"87",
   197 => x"ff",
   198 => x"c0",
   199 => x"87",
   200 => x"0e",
   201 => x"5e",
   202 => x"5b",
   203 => x"5c",
   204 => x"5d",
   205 => x"0e",
   206 => x"f0",
   207 => x"86",
   208 => x"c7",
   209 => x"ff",
   210 => x"49",
   211 => x"c0",
   212 => x"f3",
   213 => x"e1",
   214 => x"87",
   215 => x"d2",
   216 => x"c3",
   217 => x"87",
   218 => x"70",
   219 => x"98",
   220 => x"02",
   221 => x"c3",
   222 => x"cc",
   223 => x"87",
   224 => x"c7",
   225 => x"e8",
   226 => x"49",
   227 => x"c0",
   228 => x"f3",
   229 => x"d1",
   230 => x"87",
   231 => x"d8",
   232 => x"d2",
   233 => x"87",
   234 => x"70",
   235 => x"98",
   236 => x"02",
   237 => x"c2",
   238 => x"f5",
   239 => x"87",
   240 => x"c2",
   241 => x"c0",
   242 => x"c0",
   243 => x"1e",
   244 => x"c7",
   245 => x"c0",
   246 => x"49",
   247 => x"c0",
   248 => x"f0",
   249 => x"c6",
   250 => x"87",
   251 => x"c4",
   252 => x"86",
   253 => x"70",
   254 => x"4b",
   255 => x"73",
   256 => x"9b",
   257 => x"02",
   258 => x"c2",
   259 => x"e7",
   260 => x"87",
   261 => x"c4",
   262 => x"a6",
   263 => x"48",
   264 => x"c0",
   265 => x"78",
   266 => x"c4",
   267 => x"80",
   268 => x"c2",
   269 => x"c0",
   270 => x"c0",
   271 => x"78",
   272 => x"c0",
   273 => x"4d",
   274 => x"c3",
   275 => x"83",
   276 => x"fc",
   277 => x"9b",
   278 => x"c2",
   279 => x"c0",
   280 => x"c0",
   281 => x"4c",
   282 => x"73",
   283 => x"84",
   284 => x"74",
   285 => x"1e",
   286 => x"c6",
   287 => x"f4",
   288 => x"49",
   289 => x"c0",
   290 => x"ef",
   291 => x"dc",
   292 => x"87",
   293 => x"c4",
   294 => x"86",
   295 => x"70",
   296 => x"98",
   297 => x"02",
   298 => x"c1",
   299 => x"ed",
   300 => x"87",
   301 => x"c7",
   302 => x"ff",
   303 => x"b7",
   304 => x"ab",
   305 => x"06",
   306 => x"c1",
   307 => x"e5",
   308 => x"87",
   309 => x"c8",
   310 => x"c0",
   311 => x"1e",
   312 => x"cc",
   313 => x"66",
   314 => x"49",
   315 => x"75",
   316 => x"81",
   317 => x"c0",
   318 => x"f2",
   319 => x"e1",
   320 => x"87",
   321 => x"c4",
   322 => x"86",
   323 => x"70",
   324 => x"49",
   325 => x"d0",
   326 => x"a6",
   327 => x"59",
   328 => x"24",
   329 => x"7e",
   330 => x"c8",
   331 => x"c0",
   332 => x"85",
   333 => x"8b",
   334 => x"cc",
   335 => x"66",
   336 => x"48",
   337 => x"6e",
   338 => x"a8",
   339 => x"02",
   340 => x"c0",
   341 => x"fb",
   342 => x"87",
   343 => x"c4",
   344 => x"66",
   345 => x"48",
   346 => x"c1",
   347 => x"80",
   348 => x"c8",
   349 => x"a6",
   350 => x"58",
   351 => x"c1",
   352 => x"c7",
   353 => x"e8",
   354 => x"1e",
   355 => x"75",
   356 => x"49",
   357 => x"fc",
   358 => x"e6",
   359 => x"87",
   360 => x"c1",
   361 => x"c7",
   362 => x"f0",
   363 => x"48",
   364 => x"c0",
   365 => x"e0",
   366 => x"50",
   367 => x"c1",
   368 => x"c7",
   369 => x"f1",
   370 => x"1e",
   371 => x"d4",
   372 => x"66",
   373 => x"49",
   374 => x"fc",
   375 => x"d5",
   376 => x"87",
   377 => x"c1",
   378 => x"c7",
   379 => x"f9",
   380 => x"48",
   381 => x"c0",
   382 => x"e0",
   383 => x"50",
   384 => x"c1",
   385 => x"c7",
   386 => x"fa",
   387 => x"1e",
   388 => x"cc",
   389 => x"66",
   390 => x"49",
   391 => x"fc",
   392 => x"c4",
   393 => x"87",
   394 => x"cc",
   395 => x"86",
   396 => x"c1",
   397 => x"c8",
   398 => x"c2",
   399 => x"48",
   400 => x"c0",
   401 => x"50",
   402 => x"c7",
   403 => x"ff",
   404 => x"b7",
   405 => x"ab",
   406 => x"01",
   407 => x"fe",
   408 => x"db",
   409 => x"87",
   410 => x"c4",
   411 => x"66",
   412 => x"05",
   413 => x"cd",
   414 => x"87",
   415 => x"fb",
   416 => x"d9",
   417 => x"87",
   418 => x"c0",
   419 => x"c7",
   420 => x"87",
   421 => x"c7",
   422 => x"cc",
   423 => x"49",
   424 => x"c0",
   425 => x"f0",
   426 => x"cc",
   427 => x"87",
   428 => x"ff",
   429 => x"fd",
   430 => x"87",
   431 => x"f0",
   432 => x"8e",
   433 => x"fb",
   434 => x"d2",
   435 => x"87",
   436 => x"43",
   437 => x"48",
   438 => x"45",
   439 => x"43",
   440 => x"4b",
   441 => x"53",
   442 => x"55",
   443 => x"4d",
   444 => x"42",
   445 => x"49",
   446 => x"4e",
   447 => x"00",
   448 => x"38",
   449 => x"33",
   450 => x"32",
   451 => x"4f",
   452 => x"53",
   453 => x"44",
   454 => x"41",
   455 => x"41",
   456 => x"42",
   457 => x"49",
   458 => x"4e",
   459 => x"00",
   460 => x"55",
   461 => x"6e",
   462 => x"61",
   463 => x"62",
   464 => x"6c",
   465 => x"65",
   466 => x"20",
   467 => x"74",
   468 => x"6f",
   469 => x"20",
   470 => x"6c",
   471 => x"6f",
   472 => x"63",
   473 => x"61",
   474 => x"74",
   475 => x"65",
   476 => x"20",
   477 => x"70",
   478 => x"61",
   479 => x"72",
   480 => x"74",
   481 => x"69",
   482 => x"74",
   483 => x"69",
   484 => x"6f",
   485 => x"6e",
   486 => x"0a",
   487 => x"00",
   488 => x"48",
   489 => x"75",
   490 => x"6e",
   491 => x"74",
   492 => x"69",
   493 => x"6e",
   494 => x"67",
   495 => x"20",
   496 => x"66",
   497 => x"6f",
   498 => x"72",
   499 => x"20",
   500 => x"70",
   501 => x"61",
   502 => x"72",
   503 => x"74",
   504 => x"69",
   505 => x"74",
   506 => x"69",
   507 => x"6f",
   508 => x"6e",
   509 => x"0a",
   510 => x"00",
   511 => x"49",
   512 => x"6e",
   513 => x"69",
   514 => x"74",
   515 => x"69",
   516 => x"61",
   517 => x"6c",
   518 => x"69",
   519 => x"7a",
   520 => x"69",
   521 => x"6e",
   522 => x"67",
   523 => x"20",
   524 => x"53",
   525 => x"44",
   526 => x"20",
   527 => x"63",
   528 => x"61",
   529 => x"72",
   530 => x"64",
   531 => x"0a",
   532 => x"00",
   533 => x"1e",
   534 => x"e4",
   535 => x"86",
   536 => x"c0",
   537 => x"f6",
   538 => x"e4",
   539 => x"c0",
   540 => x"c0",
   541 => x"4a",
   542 => x"c3",
   543 => x"ff",
   544 => x"97",
   545 => x"7a",
   546 => x"97",
   547 => x"6a",
   548 => x"48",
   549 => x"c4",
   550 => x"a6",
   551 => x"58",
   552 => x"6e",
   553 => x"49",
   554 => x"c3",
   555 => x"ff",
   556 => x"99",
   557 => x"97",
   558 => x"7a",
   559 => x"c8",
   560 => x"31",
   561 => x"97",
   562 => x"6a",
   563 => x"48",
   564 => x"c8",
   565 => x"a6",
   566 => x"58",
   567 => x"c4",
   568 => x"66",
   569 => x"48",
   570 => x"c3",
   571 => x"ff",
   572 => x"98",
   573 => x"cc",
   574 => x"a6",
   575 => x"58",
   576 => x"c8",
   577 => x"66",
   578 => x"b1",
   579 => x"c3",
   580 => x"ff",
   581 => x"97",
   582 => x"7a",
   583 => x"c8",
   584 => x"31",
   585 => x"97",
   586 => x"6a",
   587 => x"48",
   588 => x"d0",
   589 => x"a6",
   590 => x"58",
   591 => x"cc",
   592 => x"66",
   593 => x"48",
   594 => x"c3",
   595 => x"ff",
   596 => x"98",
   597 => x"d4",
   598 => x"a6",
   599 => x"58",
   600 => x"d0",
   601 => x"66",
   602 => x"b1",
   603 => x"c3",
   604 => x"ff",
   605 => x"97",
   606 => x"7a",
   607 => x"c8",
   608 => x"31",
   609 => x"12",
   610 => x"48",
   611 => x"d8",
   612 => x"a6",
   613 => x"58",
   614 => x"d4",
   615 => x"66",
   616 => x"48",
   617 => x"c3",
   618 => x"ff",
   619 => x"98",
   620 => x"dc",
   621 => x"a6",
   622 => x"58",
   623 => x"d8",
   624 => x"66",
   625 => x"b1",
   626 => x"71",
   627 => x"48",
   628 => x"e4",
   629 => x"8e",
   630 => x"26",
   631 => x"4f",
   632 => x"0e",
   633 => x"5e",
   634 => x"5b",
   635 => x"5c",
   636 => x"5d",
   637 => x"0e",
   638 => x"1e",
   639 => x"71",
   640 => x"4a",
   641 => x"c0",
   642 => x"f6",
   643 => x"e4",
   644 => x"c0",
   645 => x"c0",
   646 => x"4b",
   647 => x"72",
   648 => x"49",
   649 => x"c3",
   650 => x"ff",
   651 => x"99",
   652 => x"73",
   653 => x"09",
   654 => x"97",
   655 => x"79",
   656 => x"09",
   657 => x"c1",
   658 => x"c8",
   659 => x"c8",
   660 => x"bf",
   661 => x"05",
   662 => x"c8",
   663 => x"87",
   664 => x"d4",
   665 => x"66",
   666 => x"48",
   667 => x"c9",
   668 => x"30",
   669 => x"d8",
   670 => x"a6",
   671 => x"58",
   672 => x"d4",
   673 => x"66",
   674 => x"49",
   675 => x"d8",
   676 => x"29",
   677 => x"c3",
   678 => x"ff",
   679 => x"99",
   680 => x"73",
   681 => x"09",
   682 => x"97",
   683 => x"79",
   684 => x"09",
   685 => x"d4",
   686 => x"66",
   687 => x"49",
   688 => x"d0",
   689 => x"29",
   690 => x"c3",
   691 => x"ff",
   692 => x"99",
   693 => x"73",
   694 => x"09",
   695 => x"97",
   696 => x"79",
   697 => x"09",
   698 => x"d4",
   699 => x"66",
   700 => x"49",
   701 => x"c8",
   702 => x"29",
   703 => x"c3",
   704 => x"ff",
   705 => x"99",
   706 => x"73",
   707 => x"09",
   708 => x"97",
   709 => x"79",
   710 => x"09",
   711 => x"d4",
   712 => x"66",
   713 => x"49",
   714 => x"c3",
   715 => x"ff",
   716 => x"99",
   717 => x"73",
   718 => x"09",
   719 => x"97",
   720 => x"79",
   721 => x"09",
   722 => x"72",
   723 => x"49",
   724 => x"d0",
   725 => x"29",
   726 => x"c3",
   727 => x"ff",
   728 => x"99",
   729 => x"73",
   730 => x"09",
   731 => x"97",
   732 => x"79",
   733 => x"09",
   734 => x"97",
   735 => x"6b",
   736 => x"48",
   737 => x"c4",
   738 => x"a6",
   739 => x"58",
   740 => x"6e",
   741 => x"4c",
   742 => x"c3",
   743 => x"ff",
   744 => x"9c",
   745 => x"c9",
   746 => x"f0",
   747 => x"ff",
   748 => x"4d",
   749 => x"c3",
   750 => x"ff",
   751 => x"ac",
   752 => x"05",
   753 => x"da",
   754 => x"87",
   755 => x"c3",
   756 => x"ff",
   757 => x"97",
   758 => x"7b",
   759 => x"97",
   760 => x"6b",
   761 => x"48",
   762 => x"c4",
   763 => x"a6",
   764 => x"58",
   765 => x"6e",
   766 => x"4c",
   767 => x"c3",
   768 => x"ff",
   769 => x"9c",
   770 => x"c1",
   771 => x"8d",
   772 => x"02",
   773 => x"c6",
   774 => x"87",
   775 => x"c3",
   776 => x"ff",
   777 => x"ac",
   778 => x"02",
   779 => x"e6",
   780 => x"87",
   781 => x"74",
   782 => x"4a",
   783 => x"c4",
   784 => x"b7",
   785 => x"2a",
   786 => x"c0",
   787 => x"f0",
   788 => x"a2",
   789 => x"49",
   790 => x"c0",
   791 => x"ea",
   792 => x"d0",
   793 => x"87",
   794 => x"74",
   795 => x"4a",
   796 => x"cf",
   797 => x"9a",
   798 => x"c0",
   799 => x"f0",
   800 => x"a2",
   801 => x"49",
   802 => x"c0",
   803 => x"ea",
   804 => x"c4",
   805 => x"87",
   806 => x"74",
   807 => x"48",
   808 => x"26",
   809 => x"26",
   810 => x"4d",
   811 => x"26",
   812 => x"4c",
   813 => x"26",
   814 => x"4b",
   815 => x"26",
   816 => x"4f",
   817 => x"1e",
   818 => x"c0",
   819 => x"49",
   820 => x"c0",
   821 => x"f6",
   822 => x"e4",
   823 => x"c0",
   824 => x"c0",
   825 => x"48",
   826 => x"c3",
   827 => x"ff",
   828 => x"50",
   829 => x"c1",
   830 => x"81",
   831 => x"c3",
   832 => x"c8",
   833 => x"b7",
   834 => x"a9",
   835 => x"04",
   836 => x"ee",
   837 => x"87",
   838 => x"26",
   839 => x"4f",
   840 => x"0e",
   841 => x"5e",
   842 => x"5b",
   843 => x"5c",
   844 => x"0e",
   845 => x"c0",
   846 => x"f6",
   847 => x"e4",
   848 => x"c0",
   849 => x"c0",
   850 => x"4c",
   851 => x"ff",
   852 => x"db",
   853 => x"87",
   854 => x"c4",
   855 => x"f8",
   856 => x"df",
   857 => x"4b",
   858 => x"c0",
   859 => x"1e",
   860 => x"c0",
   861 => x"ff",
   862 => x"f0",
   863 => x"c1",
   864 => x"f7",
   865 => x"49",
   866 => x"fc",
   867 => x"d3",
   868 => x"87",
   869 => x"c4",
   870 => x"86",
   871 => x"c1",
   872 => x"a8",
   873 => x"05",
   874 => x"c0",
   875 => x"e6",
   876 => x"87",
   877 => x"c3",
   878 => x"ff",
   879 => x"97",
   880 => x"7c",
   881 => x"c1",
   882 => x"c0",
   883 => x"c0",
   884 => x"c0",
   885 => x"c0",
   886 => x"c0",
   887 => x"1e",
   888 => x"c0",
   889 => x"e1",
   890 => x"f0",
   891 => x"c1",
   892 => x"e9",
   893 => x"49",
   894 => x"fb",
   895 => x"f7",
   896 => x"87",
   897 => x"c4",
   898 => x"86",
   899 => x"70",
   900 => x"98",
   901 => x"05",
   902 => x"c8",
   903 => x"87",
   904 => x"c3",
   905 => x"ff",
   906 => x"97",
   907 => x"7c",
   908 => x"c1",
   909 => x"48",
   910 => x"cb",
   911 => x"87",
   912 => x"fe",
   913 => x"de",
   914 => x"87",
   915 => x"c1",
   916 => x"8b",
   917 => x"05",
   918 => x"ff",
   919 => x"c1",
   920 => x"87",
   921 => x"c0",
   922 => x"48",
   923 => x"fe",
   924 => x"cd",
   925 => x"87",
   926 => x"43",
   927 => x"4d",
   928 => x"44",
   929 => x"34",
   930 => x"31",
   931 => x"20",
   932 => x"25",
   933 => x"64",
   934 => x"0a",
   935 => x"00",
   936 => x"43",
   937 => x"4d",
   938 => x"44",
   939 => x"35",
   940 => x"35",
   941 => x"20",
   942 => x"25",
   943 => x"64",
   944 => x"0a",
   945 => x"00",
   946 => x"43",
   947 => x"4d",
   948 => x"44",
   949 => x"34",
   950 => x"31",
   951 => x"20",
   952 => x"25",
   953 => x"64",
   954 => x"0a",
   955 => x"00",
   956 => x"43",
   957 => x"4d",
   958 => x"44",
   959 => x"35",
   960 => x"35",
   961 => x"20",
   962 => x"25",
   963 => x"64",
   964 => x"0a",
   965 => x"00",
   966 => x"69",
   967 => x"6e",
   968 => x"69",
   969 => x"74",
   970 => x"20",
   971 => x"25",
   972 => x"64",
   973 => x"0a",
   974 => x"20",
   975 => x"20",
   976 => x"00",
   977 => x"69",
   978 => x"6e",
   979 => x"69",
   980 => x"74",
   981 => x"20",
   982 => x"25",
   983 => x"64",
   984 => x"0a",
   985 => x"20",
   986 => x"20",
   987 => x"00",
   988 => x"43",
   989 => x"6d",
   990 => x"64",
   991 => x"5f",
   992 => x"69",
   993 => x"6e",
   994 => x"69",
   995 => x"74",
   996 => x"0a",
   997 => x"00",
   998 => x"43",
   999 => x"4d",
  1000 => x"44",
  1001 => x"38",
  1002 => x"5f",
  1003 => x"34",
  1004 => x"20",
  1005 => x"72",
  1006 => x"65",
  1007 => x"73",
  1008 => x"70",
  1009 => x"6f",
  1010 => x"6e",
  1011 => x"73",
  1012 => x"65",
  1013 => x"3a",
  1014 => x"20",
  1015 => x"25",
  1016 => x"64",
  1017 => x"0a",
  1018 => x"00",
  1019 => x"43",
  1020 => x"4d",
  1021 => x"44",
  1022 => x"35",
  1023 => x"38",
  1024 => x"20",
  1025 => x"25",
  1026 => x"64",
  1027 => x"0a",
  1028 => x"20",
  1029 => x"20",
  1030 => x"00",
  1031 => x"43",
  1032 => x"4d",
  1033 => x"44",
  1034 => x"35",
  1035 => x"38",
  1036 => x"5f",
  1037 => x"32",
  1038 => x"20",
  1039 => x"25",
  1040 => x"64",
  1041 => x"0a",
  1042 => x"20",
  1043 => x"20",
  1044 => x"00",
  1045 => x"43",
  1046 => x"4d",
  1047 => x"44",
  1048 => x"35",
  1049 => x"38",
  1050 => x"20",
  1051 => x"25",
  1052 => x"64",
  1053 => x"0a",
  1054 => x"20",
  1055 => x"20",
  1056 => x"00",
  1057 => x"53",
  1058 => x"44",
  1059 => x"48",
  1060 => x"43",
  1061 => x"20",
  1062 => x"49",
  1063 => x"6e",
  1064 => x"69",
  1065 => x"74",
  1066 => x"69",
  1067 => x"61",
  1068 => x"6c",
  1069 => x"69",
  1070 => x"7a",
  1071 => x"61",
  1072 => x"74",
  1073 => x"69",
  1074 => x"6f",
  1075 => x"6e",
  1076 => x"20",
  1077 => x"65",
  1078 => x"72",
  1079 => x"72",
  1080 => x"6f",
  1081 => x"72",
  1082 => x"21",
  1083 => x"0a",
  1084 => x"00",
  1085 => x"63",
  1086 => x"6d",
  1087 => x"64",
  1088 => x"5f",
  1089 => x"43",
  1090 => x"4d",
  1091 => x"44",
  1092 => x"38",
  1093 => x"20",
  1094 => x"72",
  1095 => x"65",
  1096 => x"73",
  1097 => x"70",
  1098 => x"6f",
  1099 => x"6e",
  1100 => x"73",
  1101 => x"65",
  1102 => x"3a",
  1103 => x"20",
  1104 => x"25",
  1105 => x"64",
  1106 => x"0a",
  1107 => x"00",
  1108 => x"52",
  1109 => x"65",
  1110 => x"61",
  1111 => x"64",
  1112 => x"20",
  1113 => x"63",
  1114 => x"6f",
  1115 => x"6d",
  1116 => x"6d",
  1117 => x"61",
  1118 => x"6e",
  1119 => x"64",
  1120 => x"20",
  1121 => x"66",
  1122 => x"61",
  1123 => x"69",
  1124 => x"6c",
  1125 => x"65",
  1126 => x"64",
  1127 => x"20",
  1128 => x"61",
  1129 => x"74",
  1130 => x"20",
  1131 => x"25",
  1132 => x"64",
  1133 => x"20",
  1134 => x"28",
  1135 => x"25",
  1136 => x"64",
  1137 => x"29",
  1138 => x"0a",
  1139 => x"00",
  1140 => x"0e",
  1141 => x"5e",
  1142 => x"5b",
  1143 => x"5c",
  1144 => x"0e",
  1145 => x"c0",
  1146 => x"f6",
  1147 => x"e4",
  1148 => x"c0",
  1149 => x"c0",
  1150 => x"4c",
  1151 => x"c3",
  1152 => x"ff",
  1153 => x"97",
  1154 => x"7c",
  1155 => x"cf",
  1156 => x"dc",
  1157 => x"49",
  1158 => x"c0",
  1159 => x"e4",
  1160 => x"ee",
  1161 => x"87",
  1162 => x"d3",
  1163 => x"4b",
  1164 => x"c0",
  1165 => x"1e",
  1166 => x"c0",
  1167 => x"ff",
  1168 => x"f0",
  1169 => x"c1",
  1170 => x"c1",
  1171 => x"49",
  1172 => x"f7",
  1173 => x"e1",
  1174 => x"87",
  1175 => x"c4",
  1176 => x"86",
  1177 => x"70",
  1178 => x"98",
  1179 => x"05",
  1180 => x"c8",
  1181 => x"87",
  1182 => x"c3",
  1183 => x"ff",
  1184 => x"97",
  1185 => x"7c",
  1186 => x"c1",
  1187 => x"48",
  1188 => x"cb",
  1189 => x"87",
  1190 => x"fa",
  1191 => x"c8",
  1192 => x"87",
  1193 => x"c1",
  1194 => x"8b",
  1195 => x"05",
  1196 => x"ff",
  1197 => x"dd",
  1198 => x"87",
  1199 => x"c0",
  1200 => x"48",
  1201 => x"f9",
  1202 => x"f7",
  1203 => x"87",
  1204 => x"0e",
  1205 => x"5e",
  1206 => x"5b",
  1207 => x"5c",
  1208 => x"0e",
  1209 => x"1e",
  1210 => x"c0",
  1211 => x"f6",
  1212 => x"e4",
  1213 => x"c0",
  1214 => x"c0",
  1215 => x"4c",
  1216 => x"f9",
  1217 => x"ee",
  1218 => x"87",
  1219 => x"c6",
  1220 => x"ea",
  1221 => x"1e",
  1222 => x"c0",
  1223 => x"e1",
  1224 => x"f0",
  1225 => x"c1",
  1226 => x"c8",
  1227 => x"49",
  1228 => x"f6",
  1229 => x"e9",
  1230 => x"87",
  1231 => x"70",
  1232 => x"4b",
  1233 => x"73",
  1234 => x"1e",
  1235 => x"d0",
  1236 => x"fd",
  1237 => x"49",
  1238 => x"c0",
  1239 => x"f2",
  1240 => x"d5",
  1241 => x"87",
  1242 => x"c8",
  1243 => x"86",
  1244 => x"c1",
  1245 => x"ab",
  1246 => x"02",
  1247 => x"c8",
  1248 => x"87",
  1249 => x"fe",
  1250 => x"d0",
  1251 => x"87",
  1252 => x"c0",
  1253 => x"48",
  1254 => x"c1",
  1255 => x"f0",
  1256 => x"87",
  1257 => x"f4",
  1258 => x"e9",
  1259 => x"87",
  1260 => x"70",
  1261 => x"49",
  1262 => x"cf",
  1263 => x"ff",
  1264 => x"ff",
  1265 => x"99",
  1266 => x"c6",
  1267 => x"ea",
  1268 => x"a9",
  1269 => x"02",
  1270 => x"c8",
  1271 => x"87",
  1272 => x"fd",
  1273 => x"f9",
  1274 => x"87",
  1275 => x"c0",
  1276 => x"48",
  1277 => x"c1",
  1278 => x"d9",
  1279 => x"87",
  1280 => x"c3",
  1281 => x"ff",
  1282 => x"97",
  1283 => x"7c",
  1284 => x"c0",
  1285 => x"f1",
  1286 => x"4b",
  1287 => x"f8",
  1288 => x"fe",
  1289 => x"87",
  1290 => x"70",
  1291 => x"98",
  1292 => x"02",
  1293 => x"c0",
  1294 => x"f8",
  1295 => x"87",
  1296 => x"c0",
  1297 => x"1e",
  1298 => x"c0",
  1299 => x"ff",
  1300 => x"f0",
  1301 => x"c1",
  1302 => x"fa",
  1303 => x"49",
  1304 => x"f5",
  1305 => x"dd",
  1306 => x"87",
  1307 => x"c4",
  1308 => x"86",
  1309 => x"70",
  1310 => x"98",
  1311 => x"05",
  1312 => x"c0",
  1313 => x"e5",
  1314 => x"87",
  1315 => x"c3",
  1316 => x"ff",
  1317 => x"97",
  1318 => x"7c",
  1319 => x"97",
  1320 => x"6c",
  1321 => x"48",
  1322 => x"c4",
  1323 => x"a6",
  1324 => x"58",
  1325 => x"6e",
  1326 => x"49",
  1327 => x"c3",
  1328 => x"ff",
  1329 => x"99",
  1330 => x"97",
  1331 => x"7c",
  1332 => x"97",
  1333 => x"7c",
  1334 => x"97",
  1335 => x"7c",
  1336 => x"97",
  1337 => x"7c",
  1338 => x"c1",
  1339 => x"c0",
  1340 => x"99",
  1341 => x"02",
  1342 => x"c4",
  1343 => x"87",
  1344 => x"c1",
  1345 => x"48",
  1346 => x"d5",
  1347 => x"87",
  1348 => x"c0",
  1349 => x"48",
  1350 => x"d1",
  1351 => x"87",
  1352 => x"c2",
  1353 => x"ab",
  1354 => x"05",
  1355 => x"c4",
  1356 => x"87",
  1357 => x"c0",
  1358 => x"48",
  1359 => x"c8",
  1360 => x"87",
  1361 => x"c1",
  1362 => x"8b",
  1363 => x"05",
  1364 => x"fe",
  1365 => x"f0",
  1366 => x"87",
  1367 => x"c0",
  1368 => x"48",
  1369 => x"26",
  1370 => x"f7",
  1371 => x"ce",
  1372 => x"87",
  1373 => x"0e",
  1374 => x"5e",
  1375 => x"5b",
  1376 => x"5c",
  1377 => x"5d",
  1378 => x"0e",
  1379 => x"c0",
  1380 => x"f6",
  1381 => x"e4",
  1382 => x"c0",
  1383 => x"c0",
  1384 => x"4c",
  1385 => x"48",
  1386 => x"c4",
  1387 => x"a0",
  1388 => x"4b",
  1389 => x"c1",
  1390 => x"c8",
  1391 => x"c8",
  1392 => x"48",
  1393 => x"c1",
  1394 => x"78",
  1395 => x"c0",
  1396 => x"f6",
  1397 => x"e4",
  1398 => x"c0",
  1399 => x"c8",
  1400 => x"48",
  1401 => x"c3",
  1402 => x"ef",
  1403 => x"50",
  1404 => x"c7",
  1405 => x"4d",
  1406 => x"c3",
  1407 => x"97",
  1408 => x"7b",
  1409 => x"f6",
  1410 => x"ed",
  1411 => x"87",
  1412 => x"c2",
  1413 => x"97",
  1414 => x"7b",
  1415 => x"c3",
  1416 => x"ff",
  1417 => x"97",
  1418 => x"7c",
  1419 => x"c0",
  1420 => x"1e",
  1421 => x"c0",
  1422 => x"e5",
  1423 => x"d0",
  1424 => x"c1",
  1425 => x"c0",
  1426 => x"49",
  1427 => x"f3",
  1428 => x"e2",
  1429 => x"87",
  1430 => x"c4",
  1431 => x"86",
  1432 => x"c1",
  1433 => x"a8",
  1434 => x"05",
  1435 => x"c2",
  1436 => x"87",
  1437 => x"c1",
  1438 => x"4d",
  1439 => x"c2",
  1440 => x"ad",
  1441 => x"05",
  1442 => x"c5",
  1443 => x"87",
  1444 => x"c0",
  1445 => x"48",
  1446 => x"c0",
  1447 => x"ec",
  1448 => x"87",
  1449 => x"c1",
  1450 => x"8d",
  1451 => x"05",
  1452 => x"ff",
  1453 => x"cf",
  1454 => x"87",
  1455 => x"fc",
  1456 => x"c2",
  1457 => x"87",
  1458 => x"c1",
  1459 => x"c8",
  1460 => x"cc",
  1461 => x"58",
  1462 => x"c1",
  1463 => x"c8",
  1464 => x"c8",
  1465 => x"bf",
  1466 => x"05",
  1467 => x"cd",
  1468 => x"87",
  1469 => x"c1",
  1470 => x"1e",
  1471 => x"c0",
  1472 => x"ff",
  1473 => x"f0",
  1474 => x"c1",
  1475 => x"d0",
  1476 => x"49",
  1477 => x"f2",
  1478 => x"f0",
  1479 => x"87",
  1480 => x"c4",
  1481 => x"86",
  1482 => x"c3",
  1483 => x"ff",
  1484 => x"97",
  1485 => x"7c",
  1486 => x"c3",
  1487 => x"53",
  1488 => x"c3",
  1489 => x"ff",
  1490 => x"54",
  1491 => x"c1",
  1492 => x"48",
  1493 => x"f5",
  1494 => x"d1",
  1495 => x"87",
  1496 => x"0e",
  1497 => x"5e",
  1498 => x"5b",
  1499 => x"5c",
  1500 => x"5d",
  1501 => x"0e",
  1502 => x"f8",
  1503 => x"86",
  1504 => x"71",
  1505 => x"4a",
  1506 => x"c0",
  1507 => x"f6",
  1508 => x"e4",
  1509 => x"c0",
  1510 => x"c0",
  1511 => x"4b",
  1512 => x"c0",
  1513 => x"7e",
  1514 => x"c3",
  1515 => x"ff",
  1516 => x"97",
  1517 => x"7b",
  1518 => x"c0",
  1519 => x"f6",
  1520 => x"e4",
  1521 => x"c0",
  1522 => x"c4",
  1523 => x"48",
  1524 => x"c2",
  1525 => x"50",
  1526 => x"c0",
  1527 => x"f6",
  1528 => x"e4",
  1529 => x"c0",
  1530 => x"c8",
  1531 => x"48",
  1532 => x"c7",
  1533 => x"50",
  1534 => x"c3",
  1535 => x"ff",
  1536 => x"97",
  1537 => x"7b",
  1538 => x"72",
  1539 => x"1e",
  1540 => x"c0",
  1541 => x"ff",
  1542 => x"f0",
  1543 => x"c1",
  1544 => x"d1",
  1545 => x"49",
  1546 => x"f1",
  1547 => x"eb",
  1548 => x"87",
  1549 => x"c4",
  1550 => x"86",
  1551 => x"70",
  1552 => x"98",
  1553 => x"05",
  1554 => x"c1",
  1555 => x"ca",
  1556 => x"87",
  1557 => x"c5",
  1558 => x"ee",
  1559 => x"cd",
  1560 => x"df",
  1561 => x"4c",
  1562 => x"c3",
  1563 => x"ff",
  1564 => x"97",
  1565 => x"7b",
  1566 => x"97",
  1567 => x"6b",
  1568 => x"48",
  1569 => x"c8",
  1570 => x"a6",
  1571 => x"58",
  1572 => x"c4",
  1573 => x"66",
  1574 => x"49",
  1575 => x"c3",
  1576 => x"ff",
  1577 => x"99",
  1578 => x"c3",
  1579 => x"fe",
  1580 => x"a9",
  1581 => x"05",
  1582 => x"de",
  1583 => x"87",
  1584 => x"c0",
  1585 => x"4d",
  1586 => x"ef",
  1587 => x"e0",
  1588 => x"87",
  1589 => x"d8",
  1590 => x"66",
  1591 => x"08",
  1592 => x"78",
  1593 => x"08",
  1594 => x"d8",
  1595 => x"66",
  1596 => x"48",
  1597 => x"c4",
  1598 => x"80",
  1599 => x"dc",
  1600 => x"a6",
  1601 => x"58",
  1602 => x"c1",
  1603 => x"85",
  1604 => x"c2",
  1605 => x"c0",
  1606 => x"b7",
  1607 => x"ad",
  1608 => x"04",
  1609 => x"e7",
  1610 => x"87",
  1611 => x"c1",
  1612 => x"4c",
  1613 => x"7e",
  1614 => x"c1",
  1615 => x"8c",
  1616 => x"05",
  1617 => x"ff",
  1618 => x"c6",
  1619 => x"87",
  1620 => x"c3",
  1621 => x"ff",
  1622 => x"53",
  1623 => x"c0",
  1624 => x"f6",
  1625 => x"e4",
  1626 => x"c0",
  1627 => x"c4",
  1628 => x"48",
  1629 => x"c3",
  1630 => x"50",
  1631 => x"6e",
  1632 => x"48",
  1633 => x"f8",
  1634 => x"8e",
  1635 => x"f3",
  1636 => x"c3",
  1637 => x"87",
  1638 => x"1e",
  1639 => x"73",
  1640 => x"1e",
  1641 => x"71",
  1642 => x"4b",
  1643 => x"73",
  1644 => x"49",
  1645 => x"d8",
  1646 => x"29",
  1647 => x"c3",
  1648 => x"ff",
  1649 => x"99",
  1650 => x"73",
  1651 => x"4a",
  1652 => x"c8",
  1653 => x"2a",
  1654 => x"cf",
  1655 => x"fc",
  1656 => x"c0",
  1657 => x"9a",
  1658 => x"72",
  1659 => x"b1",
  1660 => x"73",
  1661 => x"4a",
  1662 => x"c8",
  1663 => x"32",
  1664 => x"c0",
  1665 => x"ff",
  1666 => x"f0",
  1667 => x"c0",
  1668 => x"c0",
  1669 => x"9a",
  1670 => x"72",
  1671 => x"b1",
  1672 => x"73",
  1673 => x"4a",
  1674 => x"d8",
  1675 => x"32",
  1676 => x"ff",
  1677 => x"c0",
  1678 => x"c0",
  1679 => x"c0",
  1680 => x"c0",
  1681 => x"9a",
  1682 => x"72",
  1683 => x"b1",
  1684 => x"71",
  1685 => x"48",
  1686 => x"c4",
  1687 => x"87",
  1688 => x"26",
  1689 => x"4d",
  1690 => x"26",
  1691 => x"4c",
  1692 => x"26",
  1693 => x"4b",
  1694 => x"26",
  1695 => x"4f",
  1696 => x"1e",
  1697 => x"73",
  1698 => x"1e",
  1699 => x"71",
  1700 => x"4b",
  1701 => x"73",
  1702 => x"49",
  1703 => x"c8",
  1704 => x"29",
  1705 => x"c3",
  1706 => x"ff",
  1707 => x"99",
  1708 => x"73",
  1709 => x"4a",
  1710 => x"c8",
  1711 => x"32",
  1712 => x"cf",
  1713 => x"fc",
  1714 => x"c0",
  1715 => x"9a",
  1716 => x"72",
  1717 => x"b1",
  1718 => x"71",
  1719 => x"48",
  1720 => x"e2",
  1721 => x"87",
  1722 => x"0e",
  1723 => x"5e",
  1724 => x"5b",
  1725 => x"5c",
  1726 => x"0e",
  1727 => x"71",
  1728 => x"4b",
  1729 => x"c0",
  1730 => x"4c",
  1731 => x"d0",
  1732 => x"66",
  1733 => x"48",
  1734 => x"c0",
  1735 => x"b7",
  1736 => x"a8",
  1737 => x"06",
  1738 => x"c0",
  1739 => x"e3",
  1740 => x"87",
  1741 => x"13",
  1742 => x"4a",
  1743 => x"cc",
  1744 => x"66",
  1745 => x"97",
  1746 => x"bf",
  1747 => x"49",
  1748 => x"cc",
  1749 => x"66",
  1750 => x"48",
  1751 => x"c1",
  1752 => x"80",
  1753 => x"d0",
  1754 => x"a6",
  1755 => x"58",
  1756 => x"71",
  1757 => x"b7",
  1758 => x"aa",
  1759 => x"02",
  1760 => x"c4",
  1761 => x"87",
  1762 => x"c1",
  1763 => x"48",
  1764 => x"cc",
  1765 => x"87",
  1766 => x"c1",
  1767 => x"84",
  1768 => x"d0",
  1769 => x"66",
  1770 => x"b7",
  1771 => x"ac",
  1772 => x"04",
  1773 => x"ff",
  1774 => x"dd",
  1775 => x"87",
  1776 => x"c0",
  1777 => x"48",
  1778 => x"c2",
  1779 => x"87",
  1780 => x"26",
  1781 => x"4d",
  1782 => x"26",
  1783 => x"4c",
  1784 => x"26",
  1785 => x"4b",
  1786 => x"26",
  1787 => x"4f",
  1788 => x"0e",
  1789 => x"5e",
  1790 => x"5b",
  1791 => x"5c",
  1792 => x"5d",
  1793 => x"0e",
  1794 => x"c1",
  1795 => x"d1",
  1796 => x"ca",
  1797 => x"48",
  1798 => x"ff",
  1799 => x"78",
  1800 => x"c1",
  1801 => x"d0",
  1802 => x"da",
  1803 => x"48",
  1804 => x"c0",
  1805 => x"78",
  1806 => x"c0",
  1807 => x"e9",
  1808 => x"f1",
  1809 => x"49",
  1810 => x"da",
  1811 => x"e3",
  1812 => x"87",
  1813 => x"c1",
  1814 => x"c8",
  1815 => x"d2",
  1816 => x"1e",
  1817 => x"c0",
  1818 => x"49",
  1819 => x"fa",
  1820 => x"fa",
  1821 => x"87",
  1822 => x"c4",
  1823 => x"86",
  1824 => x"70",
  1825 => x"98",
  1826 => x"05",
  1827 => x"c5",
  1828 => x"87",
  1829 => x"c0",
  1830 => x"48",
  1831 => x"cb",
  1832 => x"c1",
  1833 => x"87",
  1834 => x"c0",
  1835 => x"4b",
  1836 => x"c1",
  1837 => x"d1",
  1838 => x"c6",
  1839 => x"48",
  1840 => x"c1",
  1841 => x"78",
  1842 => x"c8",
  1843 => x"1e",
  1844 => x"c0",
  1845 => x"e9",
  1846 => x"fe",
  1847 => x"1e",
  1848 => x"c1",
  1849 => x"c9",
  1850 => x"c8",
  1851 => x"49",
  1852 => x"fd",
  1853 => x"fb",
  1854 => x"87",
  1855 => x"c8",
  1856 => x"86",
  1857 => x"70",
  1858 => x"98",
  1859 => x"05",
  1860 => x"c6",
  1861 => x"87",
  1862 => x"c1",
  1863 => x"d1",
  1864 => x"c6",
  1865 => x"48",
  1866 => x"c0",
  1867 => x"78",
  1868 => x"c8",
  1869 => x"1e",
  1870 => x"c0",
  1871 => x"ea",
  1872 => x"c7",
  1873 => x"1e",
  1874 => x"c1",
  1875 => x"c9",
  1876 => x"e4",
  1877 => x"49",
  1878 => x"fd",
  1879 => x"e1",
  1880 => x"87",
  1881 => x"c8",
  1882 => x"86",
  1883 => x"70",
  1884 => x"98",
  1885 => x"05",
  1886 => x"c6",
  1887 => x"87",
  1888 => x"c1",
  1889 => x"d1",
  1890 => x"c6",
  1891 => x"48",
  1892 => x"c0",
  1893 => x"78",
  1894 => x"c8",
  1895 => x"1e",
  1896 => x"c0",
  1897 => x"ea",
  1898 => x"d0",
  1899 => x"1e",
  1900 => x"c1",
  1901 => x"c9",
  1902 => x"e4",
  1903 => x"49",
  1904 => x"fd",
  1905 => x"c7",
  1906 => x"87",
  1907 => x"c8",
  1908 => x"86",
  1909 => x"70",
  1910 => x"98",
  1911 => x"05",
  1912 => x"c5",
  1913 => x"87",
  1914 => x"c0",
  1915 => x"48",
  1916 => x"c9",
  1917 => x"ec",
  1918 => x"87",
  1919 => x"c1",
  1920 => x"d1",
  1921 => x"c6",
  1922 => x"bf",
  1923 => x"1e",
  1924 => x"c0",
  1925 => x"ea",
  1926 => x"d9",
  1927 => x"1e",
  1928 => x"c0",
  1929 => x"e7",
  1930 => x"e3",
  1931 => x"87",
  1932 => x"c8",
  1933 => x"86",
  1934 => x"c1",
  1935 => x"d1",
  1936 => x"c6",
  1937 => x"bf",
  1938 => x"02",
  1939 => x"c1",
  1940 => x"f4",
  1941 => x"87",
  1942 => x"c1",
  1943 => x"c8",
  1944 => x"d2",
  1945 => x"4d",
  1946 => x"48",
  1947 => x"c6",
  1948 => x"fe",
  1949 => x"a0",
  1950 => x"4c",
  1951 => x"c8",
  1952 => x"c0",
  1953 => x"1e",
  1954 => x"70",
  1955 => x"49",
  1956 => x"da",
  1957 => x"e2",
  1958 => x"87",
  1959 => x"c4",
  1960 => x"86",
  1961 => x"c8",
  1962 => x"a4",
  1963 => x"49",
  1964 => x"69",
  1965 => x"4b",
  1966 => x"c1",
  1967 => x"d0",
  1968 => x"d0",
  1969 => x"9f",
  1970 => x"bf",
  1971 => x"49",
  1972 => x"c5",
  1973 => x"d6",
  1974 => x"ea",
  1975 => x"a9",
  1976 => x"05",
  1977 => x"c0",
  1978 => x"cc",
  1979 => x"87",
  1980 => x"c8",
  1981 => x"a4",
  1982 => x"4a",
  1983 => x"6a",
  1984 => x"49",
  1985 => x"fa",
  1986 => x"e2",
  1987 => x"87",
  1988 => x"70",
  1989 => x"4b",
  1990 => x"db",
  1991 => x"87",
  1992 => x"c7",
  1993 => x"fe",
  1994 => x"a5",
  1995 => x"49",
  1996 => x"9f",
  1997 => x"69",
  1998 => x"49",
  1999 => x"ca",
  2000 => x"e9",
  2001 => x"d5",
  2002 => x"a9",
  2003 => x"02",
  2004 => x"c0",
  2005 => x"cc",
  2006 => x"87",
  2007 => x"c0",
  2008 => x"e7",
  2009 => x"ee",
  2010 => x"49",
  2011 => x"d7",
  2012 => x"da",
  2013 => x"87",
  2014 => x"c0",
  2015 => x"48",
  2016 => x"c8",
  2017 => x"c8",
  2018 => x"87",
  2019 => x"73",
  2020 => x"1e",
  2021 => x"c0",
  2022 => x"e8",
  2023 => x"cc",
  2024 => x"1e",
  2025 => x"c0",
  2026 => x"e6",
  2027 => x"c2",
  2028 => x"87",
  2029 => x"c1",
  2030 => x"c8",
  2031 => x"d2",
  2032 => x"1e",
  2033 => x"73",
  2034 => x"49",
  2035 => x"f7",
  2036 => x"e2",
  2037 => x"87",
  2038 => x"cc",
  2039 => x"86",
  2040 => x"70",
  2041 => x"98",
  2042 => x"05",
  2043 => x"c0",
  2044 => x"c5",
  2045 => x"87",
  2046 => x"c0",
  2047 => x"48",
  2048 => x"c7",
  2049 => x"e8",
  2050 => x"87",
  2051 => x"c0",
  2052 => x"e8",
  2053 => x"e4",
  2054 => x"49",
  2055 => x"d6",
  2056 => x"ee",
  2057 => x"87",
  2058 => x"c8",
  2059 => x"c0",
  2060 => x"1e",
  2061 => x"c1",
  2062 => x"c8",
  2063 => x"d2",
  2064 => x"49",
  2065 => x"d8",
  2066 => x"f5",
  2067 => x"87",
  2068 => x"c0",
  2069 => x"ea",
  2070 => x"ec",
  2071 => x"1e",
  2072 => x"c0",
  2073 => x"e5",
  2074 => x"d3",
  2075 => x"87",
  2076 => x"c8",
  2077 => x"1e",
  2078 => x"c0",
  2079 => x"eb",
  2080 => x"c4",
  2081 => x"1e",
  2082 => x"c1",
  2083 => x"c9",
  2084 => x"e4",
  2085 => x"49",
  2086 => x"fa",
  2087 => x"d1",
  2088 => x"87",
  2089 => x"d0",
  2090 => x"86",
  2091 => x"70",
  2092 => x"98",
  2093 => x"05",
  2094 => x"c0",
  2095 => x"c9",
  2096 => x"87",
  2097 => x"c1",
  2098 => x"d0",
  2099 => x"da",
  2100 => x"48",
  2101 => x"c1",
  2102 => x"78",
  2103 => x"c0",
  2104 => x"e4",
  2105 => x"87",
  2106 => x"c8",
  2107 => x"1e",
  2108 => x"c0",
  2109 => x"eb",
  2110 => x"cd",
  2111 => x"1e",
  2112 => x"c1",
  2113 => x"c9",
  2114 => x"c8",
  2115 => x"49",
  2116 => x"f9",
  2117 => x"f3",
  2118 => x"87",
  2119 => x"c8",
  2120 => x"86",
  2121 => x"70",
  2122 => x"98",
  2123 => x"02",
  2124 => x"c0",
  2125 => x"cf",
  2126 => x"87",
  2127 => x"c0",
  2128 => x"e9",
  2129 => x"cb",
  2130 => x"1e",
  2131 => x"c0",
  2132 => x"e4",
  2133 => x"d8",
  2134 => x"87",
  2135 => x"c4",
  2136 => x"86",
  2137 => x"c0",
  2138 => x"48",
  2139 => x"c6",
  2140 => x"cd",
  2141 => x"87",
  2142 => x"c1",
  2143 => x"d0",
  2144 => x"d0",
  2145 => x"97",
  2146 => x"bf",
  2147 => x"49",
  2148 => x"c1",
  2149 => x"d5",
  2150 => x"a9",
  2151 => x"05",
  2152 => x"c0",
  2153 => x"cd",
  2154 => x"87",
  2155 => x"c1",
  2156 => x"d0",
  2157 => x"d1",
  2158 => x"97",
  2159 => x"bf",
  2160 => x"49",
  2161 => x"c2",
  2162 => x"ea",
  2163 => x"a9",
  2164 => x"02",
  2165 => x"c0",
  2166 => x"c5",
  2167 => x"87",
  2168 => x"c0",
  2169 => x"48",
  2170 => x"c5",
  2171 => x"ee",
  2172 => x"87",
  2173 => x"c1",
  2174 => x"c8",
  2175 => x"d2",
  2176 => x"97",
  2177 => x"bf",
  2178 => x"49",
  2179 => x"c3",
  2180 => x"e9",
  2181 => x"a9",
  2182 => x"02",
  2183 => x"c0",
  2184 => x"d2",
  2185 => x"87",
  2186 => x"c1",
  2187 => x"c8",
  2188 => x"d2",
  2189 => x"97",
  2190 => x"bf",
  2191 => x"49",
  2192 => x"c3",
  2193 => x"eb",
  2194 => x"a9",
  2195 => x"02",
  2196 => x"c0",
  2197 => x"c5",
  2198 => x"87",
  2199 => x"c0",
  2200 => x"48",
  2201 => x"c5",
  2202 => x"cf",
  2203 => x"87",
  2204 => x"c1",
  2205 => x"c8",
  2206 => x"dd",
  2207 => x"97",
  2208 => x"bf",
  2209 => x"49",
  2210 => x"71",
  2211 => x"99",
  2212 => x"05",
  2213 => x"c0",
  2214 => x"cc",
  2215 => x"87",
  2216 => x"c1",
  2217 => x"c8",
  2218 => x"de",
  2219 => x"97",
  2220 => x"bf",
  2221 => x"49",
  2222 => x"c2",
  2223 => x"a9",
  2224 => x"02",
  2225 => x"c0",
  2226 => x"c5",
  2227 => x"87",
  2228 => x"c0",
  2229 => x"48",
  2230 => x"c4",
  2231 => x"f2",
  2232 => x"87",
  2233 => x"c1",
  2234 => x"c8",
  2235 => x"df",
  2236 => x"97",
  2237 => x"bf",
  2238 => x"48",
  2239 => x"c1",
  2240 => x"d0",
  2241 => x"d6",
  2242 => x"58",
  2243 => x"c1",
  2244 => x"d0",
  2245 => x"d2",
  2246 => x"bf",
  2247 => x"48",
  2248 => x"c1",
  2249 => x"88",
  2250 => x"c1",
  2251 => x"d0",
  2252 => x"da",
  2253 => x"58",
  2254 => x"c1",
  2255 => x"c8",
  2256 => x"e0",
  2257 => x"97",
  2258 => x"bf",
  2259 => x"49",
  2260 => x"73",
  2261 => x"81",
  2262 => x"c1",
  2263 => x"c8",
  2264 => x"e1",
  2265 => x"97",
  2266 => x"bf",
  2267 => x"4a",
  2268 => x"c8",
  2269 => x"32",
  2270 => x"c1",
  2271 => x"d0",
  2272 => x"e6",
  2273 => x"48",
  2274 => x"72",
  2275 => x"a1",
  2276 => x"78",
  2277 => x"c1",
  2278 => x"c8",
  2279 => x"e2",
  2280 => x"97",
  2281 => x"bf",
  2282 => x"48",
  2283 => x"c1",
  2284 => x"d0",
  2285 => x"fe",
  2286 => x"58",
  2287 => x"c1",
  2288 => x"d0",
  2289 => x"da",
  2290 => x"bf",
  2291 => x"02",
  2292 => x"c2",
  2293 => x"e2",
  2294 => x"87",
  2295 => x"c8",
  2296 => x"1e",
  2297 => x"c0",
  2298 => x"e9",
  2299 => x"e8",
  2300 => x"1e",
  2301 => x"c1",
  2302 => x"c9",
  2303 => x"e4",
  2304 => x"49",
  2305 => x"f6",
  2306 => x"f6",
  2307 => x"87",
  2308 => x"c8",
  2309 => x"86",
  2310 => x"70",
  2311 => x"98",
  2312 => x"02",
  2313 => x"c0",
  2314 => x"c5",
  2315 => x"87",
  2316 => x"c0",
  2317 => x"48",
  2318 => x"c3",
  2319 => x"da",
  2320 => x"87",
  2321 => x"c1",
  2322 => x"d0",
  2323 => x"d2",
  2324 => x"bf",
  2325 => x"48",
  2326 => x"c4",
  2327 => x"30",
  2328 => x"c1",
  2329 => x"d1",
  2330 => x"c2",
  2331 => x"58",
  2332 => x"c1",
  2333 => x"d0",
  2334 => x"d2",
  2335 => x"bf",
  2336 => x"4a",
  2337 => x"c1",
  2338 => x"d0",
  2339 => x"fa",
  2340 => x"5a",
  2341 => x"c1",
  2342 => x"c8",
  2343 => x"f7",
  2344 => x"97",
  2345 => x"bf",
  2346 => x"49",
  2347 => x"c8",
  2348 => x"31",
  2349 => x"c1",
  2350 => x"c8",
  2351 => x"f6",
  2352 => x"97",
  2353 => x"bf",
  2354 => x"4b",
  2355 => x"73",
  2356 => x"a1",
  2357 => x"49",
  2358 => x"c1",
  2359 => x"c8",
  2360 => x"f8",
  2361 => x"97",
  2362 => x"bf",
  2363 => x"4b",
  2364 => x"d0",
  2365 => x"33",
  2366 => x"73",
  2367 => x"a1",
  2368 => x"49",
  2369 => x"c1",
  2370 => x"c8",
  2371 => x"f9",
  2372 => x"97",
  2373 => x"bf",
  2374 => x"4b",
  2375 => x"d8",
  2376 => x"33",
  2377 => x"73",
  2378 => x"a1",
  2379 => x"49",
  2380 => x"c1",
  2381 => x"d1",
  2382 => x"c6",
  2383 => x"59",
  2384 => x"c1",
  2385 => x"d0",
  2386 => x"fa",
  2387 => x"bf",
  2388 => x"91",
  2389 => x"c1",
  2390 => x"d0",
  2391 => x"e6",
  2392 => x"bf",
  2393 => x"81",
  2394 => x"c1",
  2395 => x"d0",
  2396 => x"ee",
  2397 => x"59",
  2398 => x"c1",
  2399 => x"c8",
  2400 => x"ff",
  2401 => x"97",
  2402 => x"bf",
  2403 => x"4b",
  2404 => x"c8",
  2405 => x"33",
  2406 => x"c1",
  2407 => x"c8",
  2408 => x"fe",
  2409 => x"97",
  2410 => x"bf",
  2411 => x"4c",
  2412 => x"74",
  2413 => x"a3",
  2414 => x"4b",
  2415 => x"c1",
  2416 => x"c9",
  2417 => x"c0",
  2418 => x"97",
  2419 => x"bf",
  2420 => x"4c",
  2421 => x"d0",
  2422 => x"34",
  2423 => x"74",
  2424 => x"a3",
  2425 => x"4b",
  2426 => x"c1",
  2427 => x"c9",
  2428 => x"c1",
  2429 => x"97",
  2430 => x"bf",
  2431 => x"4c",
  2432 => x"cf",
  2433 => x"9c",
  2434 => x"d8",
  2435 => x"34",
  2436 => x"74",
  2437 => x"a3",
  2438 => x"4b",
  2439 => x"c1",
  2440 => x"d0",
  2441 => x"f2",
  2442 => x"5b",
  2443 => x"c2",
  2444 => x"8b",
  2445 => x"73",
  2446 => x"92",
  2447 => x"c1",
  2448 => x"d0",
  2449 => x"f2",
  2450 => x"48",
  2451 => x"72",
  2452 => x"a1",
  2453 => x"78",
  2454 => x"c1",
  2455 => x"d0",
  2456 => x"87",
  2457 => x"c1",
  2458 => x"c8",
  2459 => x"e4",
  2460 => x"97",
  2461 => x"bf",
  2462 => x"49",
  2463 => x"c8",
  2464 => x"31",
  2465 => x"c1",
  2466 => x"c8",
  2467 => x"e3",
  2468 => x"97",
  2469 => x"bf",
  2470 => x"4a",
  2471 => x"72",
  2472 => x"a1",
  2473 => x"49",
  2474 => x"c1",
  2475 => x"d1",
  2476 => x"c2",
  2477 => x"59",
  2478 => x"c5",
  2479 => x"31",
  2480 => x"c7",
  2481 => x"ff",
  2482 => x"81",
  2483 => x"c9",
  2484 => x"29",
  2485 => x"c1",
  2486 => x"d0",
  2487 => x"fa",
  2488 => x"59",
  2489 => x"c1",
  2490 => x"c8",
  2491 => x"e9",
  2492 => x"97",
  2493 => x"bf",
  2494 => x"4a",
  2495 => x"c8",
  2496 => x"32",
  2497 => x"c1",
  2498 => x"c8",
  2499 => x"e8",
  2500 => x"97",
  2501 => x"bf",
  2502 => x"4b",
  2503 => x"73",
  2504 => x"a2",
  2505 => x"4a",
  2506 => x"c1",
  2507 => x"d1",
  2508 => x"c6",
  2509 => x"5a",
  2510 => x"c1",
  2511 => x"d0",
  2512 => x"fa",
  2513 => x"bf",
  2514 => x"92",
  2515 => x"c1",
  2516 => x"d0",
  2517 => x"e6",
  2518 => x"bf",
  2519 => x"82",
  2520 => x"c1",
  2521 => x"d0",
  2522 => x"f6",
  2523 => x"5a",
  2524 => x"c1",
  2525 => x"d0",
  2526 => x"ee",
  2527 => x"48",
  2528 => x"c0",
  2529 => x"78",
  2530 => x"c1",
  2531 => x"d0",
  2532 => x"ea",
  2533 => x"48",
  2534 => x"72",
  2535 => x"a1",
  2536 => x"78",
  2537 => x"c1",
  2538 => x"48",
  2539 => x"f4",
  2540 => x"c6",
  2541 => x"87",
  2542 => x"4e",
  2543 => x"6f",
  2544 => x"20",
  2545 => x"70",
  2546 => x"61",
  2547 => x"72",
  2548 => x"74",
  2549 => x"69",
  2550 => x"74",
  2551 => x"69",
  2552 => x"6f",
  2553 => x"6e",
  2554 => x"20",
  2555 => x"73",
  2556 => x"69",
  2557 => x"67",
  2558 => x"6e",
  2559 => x"61",
  2560 => x"74",
  2561 => x"75",
  2562 => x"72",
  2563 => x"65",
  2564 => x"20",
  2565 => x"66",
  2566 => x"6f",
  2567 => x"75",
  2568 => x"6e",
  2569 => x"64",
  2570 => x"0a",
  2571 => x"00",
  2572 => x"52",
  2573 => x"65",
  2574 => x"61",
  2575 => x"64",
  2576 => x"69",
  2577 => x"6e",
  2578 => x"67",
  2579 => x"20",
  2580 => x"62",
  2581 => x"6f",
  2582 => x"6f",
  2583 => x"74",
  2584 => x"20",
  2585 => x"73",
  2586 => x"65",
  2587 => x"63",
  2588 => x"74",
  2589 => x"6f",
  2590 => x"72",
  2591 => x"20",
  2592 => x"25",
  2593 => x"64",
  2594 => x"0a",
  2595 => x"00",
  2596 => x"52",
  2597 => x"65",
  2598 => x"61",
  2599 => x"64",
  2600 => x"20",
  2601 => x"62",
  2602 => x"6f",
  2603 => x"6f",
  2604 => x"74",
  2605 => x"20",
  2606 => x"73",
  2607 => x"65",
  2608 => x"63",
  2609 => x"74",
  2610 => x"6f",
  2611 => x"72",
  2612 => x"20",
  2613 => x"66",
  2614 => x"72",
  2615 => x"6f",
  2616 => x"6d",
  2617 => x"20",
  2618 => x"66",
  2619 => x"69",
  2620 => x"72",
  2621 => x"73",
  2622 => x"74",
  2623 => x"20",
  2624 => x"70",
  2625 => x"61",
  2626 => x"72",
  2627 => x"74",
  2628 => x"69",
  2629 => x"74",
  2630 => x"69",
  2631 => x"6f",
  2632 => x"6e",
  2633 => x"0a",
  2634 => x"00",
  2635 => x"55",
  2636 => x"6e",
  2637 => x"73",
  2638 => x"75",
  2639 => x"70",
  2640 => x"70",
  2641 => x"6f",
  2642 => x"72",
  2643 => x"74",
  2644 => x"65",
  2645 => x"64",
  2646 => x"20",
  2647 => x"70",
  2648 => x"61",
  2649 => x"72",
  2650 => x"74",
  2651 => x"69",
  2652 => x"74",
  2653 => x"69",
  2654 => x"6f",
  2655 => x"6e",
  2656 => x"20",
  2657 => x"74",
  2658 => x"79",
  2659 => x"70",
  2660 => x"65",
  2661 => x"21",
  2662 => x"0d",
  2663 => x"00",
  2664 => x"46",
  2665 => x"41",
  2666 => x"54",
  2667 => x"33",
  2668 => x"32",
  2669 => x"20",
  2670 => x"20",
  2671 => x"20",
  2672 => x"00",
  2673 => x"52",
  2674 => x"65",
  2675 => x"61",
  2676 => x"64",
  2677 => x"69",
  2678 => x"6e",
  2679 => x"67",
  2680 => x"20",
  2681 => x"4d",
  2682 => x"42",
  2683 => x"52",
  2684 => x"0a",
  2685 => x"00",
  2686 => x"46",
  2687 => x"41",
  2688 => x"54",
  2689 => x"31",
  2690 => x"36",
  2691 => x"20",
  2692 => x"20",
  2693 => x"20",
  2694 => x"00",
  2695 => x"46",
  2696 => x"41",
  2697 => x"54",
  2698 => x"33",
  2699 => x"32",
  2700 => x"20",
  2701 => x"20",
  2702 => x"20",
  2703 => x"00",
  2704 => x"46",
  2705 => x"41",
  2706 => x"54",
  2707 => x"31",
  2708 => x"32",
  2709 => x"20",
  2710 => x"20",
  2711 => x"20",
  2712 => x"00",
  2713 => x"50",
  2714 => x"61",
  2715 => x"72",
  2716 => x"74",
  2717 => x"69",
  2718 => x"74",
  2719 => x"69",
  2720 => x"6f",
  2721 => x"6e",
  2722 => x"63",
  2723 => x"6f",
  2724 => x"75",
  2725 => x"6e",
  2726 => x"74",
  2727 => x"20",
  2728 => x"25",
  2729 => x"64",
  2730 => x"0a",
  2731 => x"00",
  2732 => x"48",
  2733 => x"75",
  2734 => x"6e",
  2735 => x"74",
  2736 => x"69",
  2737 => x"6e",
  2738 => x"67",
  2739 => x"20",
  2740 => x"66",
  2741 => x"6f",
  2742 => x"72",
  2743 => x"20",
  2744 => x"66",
  2745 => x"69",
  2746 => x"6c",
  2747 => x"65",
  2748 => x"73",
  2749 => x"79",
  2750 => x"73",
  2751 => x"74",
  2752 => x"65",
  2753 => x"6d",
  2754 => x"0a",
  2755 => x"00",
  2756 => x"46",
  2757 => x"41",
  2758 => x"54",
  2759 => x"33",
  2760 => x"32",
  2761 => x"20",
  2762 => x"20",
  2763 => x"20",
  2764 => x"00",
  2765 => x"46",
  2766 => x"41",
  2767 => x"54",
  2768 => x"31",
  2769 => x"36",
  2770 => x"20",
  2771 => x"20",
  2772 => x"20",
  2773 => x"00",
  2774 => x"52",
  2775 => x"65",
  2776 => x"61",
  2777 => x"64",
  2778 => x"69",
  2779 => x"6e",
  2780 => x"67",
  2781 => x"20",
  2782 => x"64",
  2783 => x"69",
  2784 => x"72",
  2785 => x"65",
  2786 => x"63",
  2787 => x"74",
  2788 => x"6f",
  2789 => x"72",
  2790 => x"79",
  2791 => x"20",
  2792 => x"73",
  2793 => x"65",
  2794 => x"63",
  2795 => x"74",
  2796 => x"6f",
  2797 => x"72",
  2798 => x"20",
  2799 => x"25",
  2800 => x"64",
  2801 => x"0a",
  2802 => x"00",
  2803 => x"66",
  2804 => x"69",
  2805 => x"6c",
  2806 => x"65",
  2807 => x"20",
  2808 => x"22",
  2809 => x"25",
  2810 => x"73",
  2811 => x"22",
  2812 => x"20",
  2813 => x"66",
  2814 => x"6f",
  2815 => x"75",
  2816 => x"6e",
  2817 => x"64",
  2818 => x"0d",
  2819 => x"00",
  2820 => x"47",
  2821 => x"65",
  2822 => x"74",
  2823 => x"46",
  2824 => x"41",
  2825 => x"54",
  2826 => x"4c",
  2827 => x"69",
  2828 => x"6e",
  2829 => x"6b",
  2830 => x"20",
  2831 => x"72",
  2832 => x"65",
  2833 => x"74",
  2834 => x"75",
  2835 => x"72",
  2836 => x"6e",
  2837 => x"65",
  2838 => x"64",
  2839 => x"20",
  2840 => x"25",
  2841 => x"64",
  2842 => x"0a",
  2843 => x"00",
  2844 => x"43",
  2845 => x"61",
  2846 => x"6e",
  2847 => x"27",
  2848 => x"74",
  2849 => x"20",
  2850 => x"6f",
  2851 => x"70",
  2852 => x"65",
  2853 => x"6e",
  2854 => x"20",
  2855 => x"25",
  2856 => x"73",
  2857 => x"0a",
  2858 => x"00",
  2859 => x"0e",
  2860 => x"5e",
  2861 => x"5b",
  2862 => x"5c",
  2863 => x"5d",
  2864 => x"0e",
  2865 => x"71",
  2866 => x"4a",
  2867 => x"c1",
  2868 => x"d0",
  2869 => x"da",
  2870 => x"bf",
  2871 => x"02",
  2872 => x"cc",
  2873 => x"87",
  2874 => x"72",
  2875 => x"4b",
  2876 => x"c7",
  2877 => x"b7",
  2878 => x"2b",
  2879 => x"72",
  2880 => x"4c",
  2881 => x"c1",
  2882 => x"ff",
  2883 => x"9c",
  2884 => x"ca",
  2885 => x"87",
  2886 => x"72",
  2887 => x"4b",
  2888 => x"c8",
  2889 => x"b7",
  2890 => x"2b",
  2891 => x"72",
  2892 => x"4c",
  2893 => x"c3",
  2894 => x"ff",
  2895 => x"9c",
  2896 => x"c1",
  2897 => x"d1",
  2898 => x"ca",
  2899 => x"bf",
  2900 => x"ab",
  2901 => x"02",
  2902 => x"de",
  2903 => x"87",
  2904 => x"c1",
  2905 => x"c8",
  2906 => x"d2",
  2907 => x"1e",
  2908 => x"c1",
  2909 => x"d0",
  2910 => x"e6",
  2911 => x"bf",
  2912 => x"49",
  2913 => x"73",
  2914 => x"81",
  2915 => x"e9",
  2916 => x"f2",
  2917 => x"87",
  2918 => x"c4",
  2919 => x"86",
  2920 => x"70",
  2921 => x"98",
  2922 => x"05",
  2923 => x"c5",
  2924 => x"87",
  2925 => x"c0",
  2926 => x"48",
  2927 => x"c0",
  2928 => x"f6",
  2929 => x"87",
  2930 => x"c1",
  2931 => x"d1",
  2932 => x"ce",
  2933 => x"5b",
  2934 => x"c1",
  2935 => x"d0",
  2936 => x"da",
  2937 => x"bf",
  2938 => x"02",
  2939 => x"d9",
  2940 => x"87",
  2941 => x"74",
  2942 => x"4a",
  2943 => x"c4",
  2944 => x"92",
  2945 => x"c1",
  2946 => x"c8",
  2947 => x"d2",
  2948 => x"82",
  2949 => x"6a",
  2950 => x"49",
  2951 => x"eb",
  2952 => x"dc",
  2953 => x"87",
  2954 => x"70",
  2955 => x"49",
  2956 => x"71",
  2957 => x"4d",
  2958 => x"cf",
  2959 => x"ff",
  2960 => x"ff",
  2961 => x"ff",
  2962 => x"ff",
  2963 => x"9d",
  2964 => x"d0",
  2965 => x"87",
  2966 => x"74",
  2967 => x"4a",
  2968 => x"c2",
  2969 => x"92",
  2970 => x"c1",
  2971 => x"c8",
  2972 => x"d2",
  2973 => x"82",
  2974 => x"9f",
  2975 => x"6a",
  2976 => x"49",
  2977 => x"eb",
  2978 => x"fc",
  2979 => x"87",
  2980 => x"70",
  2981 => x"4d",
  2982 => x"75",
  2983 => x"48",
  2984 => x"ed",
  2985 => x"c9",
  2986 => x"87",
  2987 => x"0e",
  2988 => x"5e",
  2989 => x"5b",
  2990 => x"5c",
  2991 => x"5d",
  2992 => x"0e",
  2993 => x"f4",
  2994 => x"86",
  2995 => x"71",
  2996 => x"4c",
  2997 => x"c0",
  2998 => x"4b",
  2999 => x"c1",
  3000 => x"d1",
  3001 => x"ca",
  3002 => x"48",
  3003 => x"ff",
  3004 => x"78",
  3005 => x"c1",
  3006 => x"d0",
  3007 => x"ee",
  3008 => x"bf",
  3009 => x"4d",
  3010 => x"c1",
  3011 => x"d0",
  3012 => x"f2",
  3013 => x"bf",
  3014 => x"7e",
  3015 => x"c1",
  3016 => x"d0",
  3017 => x"da",
  3018 => x"bf",
  3019 => x"02",
  3020 => x"c9",
  3021 => x"87",
  3022 => x"c1",
  3023 => x"d0",
  3024 => x"d2",
  3025 => x"bf",
  3026 => x"4a",
  3027 => x"c4",
  3028 => x"32",
  3029 => x"c7",
  3030 => x"87",
  3031 => x"c1",
  3032 => x"d0",
  3033 => x"f6",
  3034 => x"bf",
  3035 => x"4a",
  3036 => x"c4",
  3037 => x"32",
  3038 => x"c8",
  3039 => x"a6",
  3040 => x"5a",
  3041 => x"c8",
  3042 => x"a6",
  3043 => x"48",
  3044 => x"c0",
  3045 => x"78",
  3046 => x"c4",
  3047 => x"66",
  3048 => x"48",
  3049 => x"c0",
  3050 => x"a8",
  3051 => x"06",
  3052 => x"c3",
  3053 => x"cf",
  3054 => x"87",
  3055 => x"c8",
  3056 => x"66",
  3057 => x"49",
  3058 => x"cf",
  3059 => x"99",
  3060 => x"05",
  3061 => x"c0",
  3062 => x"e3",
  3063 => x"87",
  3064 => x"6e",
  3065 => x"1e",
  3066 => x"c0",
  3067 => x"eb",
  3068 => x"d6",
  3069 => x"1e",
  3070 => x"d5",
  3071 => x"ee",
  3072 => x"87",
  3073 => x"c1",
  3074 => x"c8",
  3075 => x"d2",
  3076 => x"1e",
  3077 => x"cc",
  3078 => x"66",
  3079 => x"49",
  3080 => x"48",
  3081 => x"c1",
  3082 => x"80",
  3083 => x"d0",
  3084 => x"a6",
  3085 => x"58",
  3086 => x"71",
  3087 => x"49",
  3088 => x"e7",
  3089 => x"c5",
  3090 => x"87",
  3091 => x"cc",
  3092 => x"86",
  3093 => x"c1",
  3094 => x"c8",
  3095 => x"d2",
  3096 => x"4b",
  3097 => x"c3",
  3098 => x"87",
  3099 => x"c0",
  3100 => x"e0",
  3101 => x"83",
  3102 => x"97",
  3103 => x"6b",
  3104 => x"49",
  3105 => x"71",
  3106 => x"99",
  3107 => x"02",
  3108 => x"c2",
  3109 => x"c5",
  3110 => x"87",
  3111 => x"97",
  3112 => x"6b",
  3113 => x"49",
  3114 => x"c3",
  3115 => x"e5",
  3116 => x"a9",
  3117 => x"02",
  3118 => x"c1",
  3119 => x"fb",
  3120 => x"87",
  3121 => x"cb",
  3122 => x"a3",
  3123 => x"49",
  3124 => x"97",
  3125 => x"69",
  3126 => x"49",
  3127 => x"d8",
  3128 => x"99",
  3129 => x"05",
  3130 => x"c1",
  3131 => x"ef",
  3132 => x"87",
  3133 => x"cb",
  3134 => x"1e",
  3135 => x"c0",
  3136 => x"e0",
  3137 => x"66",
  3138 => x"1e",
  3139 => x"73",
  3140 => x"49",
  3141 => x"e9",
  3142 => x"f2",
  3143 => x"87",
  3144 => x"c8",
  3145 => x"86",
  3146 => x"70",
  3147 => x"98",
  3148 => x"05",
  3149 => x"c1",
  3150 => x"dc",
  3151 => x"87",
  3152 => x"dc",
  3153 => x"a3",
  3154 => x"4a",
  3155 => x"6a",
  3156 => x"49",
  3157 => x"e8",
  3158 => x"ce",
  3159 => x"87",
  3160 => x"70",
  3161 => x"4a",
  3162 => x"c4",
  3163 => x"a4",
  3164 => x"49",
  3165 => x"72",
  3166 => x"79",
  3167 => x"da",
  3168 => x"a3",
  3169 => x"4a",
  3170 => x"9f",
  3171 => x"6a",
  3172 => x"49",
  3173 => x"e8",
  3174 => x"f8",
  3175 => x"87",
  3176 => x"c4",
  3177 => x"a6",
  3178 => x"58",
  3179 => x"c1",
  3180 => x"d0",
  3181 => x"da",
  3182 => x"bf",
  3183 => x"02",
  3184 => x"d8",
  3185 => x"87",
  3186 => x"d4",
  3187 => x"a3",
  3188 => x"4a",
  3189 => x"9f",
  3190 => x"6a",
  3191 => x"49",
  3192 => x"e8",
  3193 => x"e5",
  3194 => x"87",
  3195 => x"70",
  3196 => x"49",
  3197 => x"c0",
  3198 => x"ff",
  3199 => x"ff",
  3200 => x"99",
  3201 => x"71",
  3202 => x"48",
  3203 => x"d0",
  3204 => x"30",
  3205 => x"c8",
  3206 => x"a6",
  3207 => x"58",
  3208 => x"c5",
  3209 => x"87",
  3210 => x"c4",
  3211 => x"a6",
  3212 => x"48",
  3213 => x"c0",
  3214 => x"78",
  3215 => x"c4",
  3216 => x"66",
  3217 => x"4a",
  3218 => x"6e",
  3219 => x"82",
  3220 => x"c8",
  3221 => x"a4",
  3222 => x"49",
  3223 => x"72",
  3224 => x"79",
  3225 => x"c0",
  3226 => x"7c",
  3227 => x"dc",
  3228 => x"66",
  3229 => x"1e",
  3230 => x"c0",
  3231 => x"eb",
  3232 => x"f3",
  3233 => x"1e",
  3234 => x"d3",
  3235 => x"ca",
  3236 => x"87",
  3237 => x"c8",
  3238 => x"86",
  3239 => x"c1",
  3240 => x"48",
  3241 => x"c1",
  3242 => x"d0",
  3243 => x"87",
  3244 => x"c8",
  3245 => x"66",
  3246 => x"48",
  3247 => x"c1",
  3248 => x"80",
  3249 => x"cc",
  3250 => x"a6",
  3251 => x"58",
  3252 => x"c8",
  3253 => x"66",
  3254 => x"48",
  3255 => x"c4",
  3256 => x"66",
  3257 => x"a8",
  3258 => x"04",
  3259 => x"fc",
  3260 => x"f1",
  3261 => x"87",
  3262 => x"c1",
  3263 => x"d0",
  3264 => x"da",
  3265 => x"bf",
  3266 => x"02",
  3267 => x"c0",
  3268 => x"f4",
  3269 => x"87",
  3270 => x"75",
  3271 => x"49",
  3272 => x"f9",
  3273 => x"e0",
  3274 => x"87",
  3275 => x"70",
  3276 => x"4d",
  3277 => x"75",
  3278 => x"1e",
  3279 => x"c0",
  3280 => x"ec",
  3281 => x"c4",
  3282 => x"1e",
  3283 => x"d2",
  3284 => x"d9",
  3285 => x"87",
  3286 => x"c8",
  3287 => x"86",
  3288 => x"75",
  3289 => x"49",
  3290 => x"cf",
  3291 => x"ff",
  3292 => x"ff",
  3293 => x"ff",
  3294 => x"f8",
  3295 => x"99",
  3296 => x"a9",
  3297 => x"02",
  3298 => x"d6",
  3299 => x"87",
  3300 => x"75",
  3301 => x"49",
  3302 => x"c2",
  3303 => x"89",
  3304 => x"c1",
  3305 => x"d0",
  3306 => x"d2",
  3307 => x"bf",
  3308 => x"91",
  3309 => x"c1",
  3310 => x"d0",
  3311 => x"ea",
  3312 => x"bf",
  3313 => x"48",
  3314 => x"71",
  3315 => x"80",
  3316 => x"c4",
  3317 => x"a6",
  3318 => x"58",
  3319 => x"fb",
  3320 => x"e7",
  3321 => x"87",
  3322 => x"c0",
  3323 => x"48",
  3324 => x"f4",
  3325 => x"8e",
  3326 => x"e7",
  3327 => x"f3",
  3328 => x"87",
  3329 => x"0e",
  3330 => x"5e",
  3331 => x"5b",
  3332 => x"5c",
  3333 => x"5d",
  3334 => x"0e",
  3335 => x"1e",
  3336 => x"71",
  3337 => x"4b",
  3338 => x"73",
  3339 => x"1e",
  3340 => x"c1",
  3341 => x"d1",
  3342 => x"ce",
  3343 => x"49",
  3344 => x"fa",
  3345 => x"d8",
  3346 => x"87",
  3347 => x"c4",
  3348 => x"86",
  3349 => x"70",
  3350 => x"98",
  3351 => x"02",
  3352 => x"c1",
  3353 => x"f7",
  3354 => x"87",
  3355 => x"c1",
  3356 => x"d1",
  3357 => x"d2",
  3358 => x"bf",
  3359 => x"49",
  3360 => x"c7",
  3361 => x"ff",
  3362 => x"81",
  3363 => x"c9",
  3364 => x"29",
  3365 => x"c4",
  3366 => x"a6",
  3367 => x"59",
  3368 => x"c0",
  3369 => x"4d",
  3370 => x"4c",
  3371 => x"6e",
  3372 => x"48",
  3373 => x"c0",
  3374 => x"b7",
  3375 => x"a8",
  3376 => x"06",
  3377 => x"c1",
  3378 => x"ed",
  3379 => x"87",
  3380 => x"c1",
  3381 => x"d0",
  3382 => x"ea",
  3383 => x"bf",
  3384 => x"49",
  3385 => x"c1",
  3386 => x"d1",
  3387 => x"d6",
  3388 => x"bf",
  3389 => x"4a",
  3390 => x"c2",
  3391 => x"8a",
  3392 => x"c1",
  3393 => x"d0",
  3394 => x"d2",
  3395 => x"bf",
  3396 => x"92",
  3397 => x"72",
  3398 => x"a1",
  3399 => x"49",
  3400 => x"c1",
  3401 => x"d0",
  3402 => x"d6",
  3403 => x"bf",
  3404 => x"4a",
  3405 => x"74",
  3406 => x"9a",
  3407 => x"72",
  3408 => x"a1",
  3409 => x"49",
  3410 => x"d4",
  3411 => x"66",
  3412 => x"1e",
  3413 => x"71",
  3414 => x"49",
  3415 => x"e1",
  3416 => x"fe",
  3417 => x"87",
  3418 => x"c4",
  3419 => x"86",
  3420 => x"70",
  3421 => x"98",
  3422 => x"05",
  3423 => x"c5",
  3424 => x"87",
  3425 => x"c0",
  3426 => x"48",
  3427 => x"c1",
  3428 => x"c0",
  3429 => x"87",
  3430 => x"c1",
  3431 => x"84",
  3432 => x"c1",
  3433 => x"d0",
  3434 => x"d6",
  3435 => x"bf",
  3436 => x"49",
  3437 => x"74",
  3438 => x"99",
  3439 => x"05",
  3440 => x"cc",
  3441 => x"87",
  3442 => x"c1",
  3443 => x"d1",
  3444 => x"d6",
  3445 => x"bf",
  3446 => x"49",
  3447 => x"f6",
  3448 => x"f1",
  3449 => x"87",
  3450 => x"c1",
  3451 => x"d1",
  3452 => x"da",
  3453 => x"58",
  3454 => x"d4",
  3455 => x"66",
  3456 => x"48",
  3457 => x"c8",
  3458 => x"c0",
  3459 => x"80",
  3460 => x"d8",
  3461 => x"a6",
  3462 => x"58",
  3463 => x"c1",
  3464 => x"85",
  3465 => x"6e",
  3466 => x"b7",
  3467 => x"ad",
  3468 => x"04",
  3469 => x"fe",
  3470 => x"e4",
  3471 => x"87",
  3472 => x"cf",
  3473 => x"87",
  3474 => x"73",
  3475 => x"1e",
  3476 => x"c0",
  3477 => x"ec",
  3478 => x"dc",
  3479 => x"1e",
  3480 => x"cf",
  3481 => x"d4",
  3482 => x"87",
  3483 => x"c8",
  3484 => x"86",
  3485 => x"c0",
  3486 => x"48",
  3487 => x"c5",
  3488 => x"87",
  3489 => x"c1",
  3490 => x"d1",
  3491 => x"d2",
  3492 => x"bf",
  3493 => x"48",
  3494 => x"26",
  3495 => x"e5",
  3496 => x"ca",
  3497 => x"87",
  3498 => x"1e",
  3499 => x"c0",
  3500 => x"f6",
  3501 => x"e8",
  3502 => x"c0",
  3503 => x"c0",
  3504 => x"09",
  3505 => x"97",
  3506 => x"79",
  3507 => x"09",
  3508 => x"71",
  3509 => x"48",
  3510 => x"26",
  3511 => x"4f",
  3512 => x"0e",
  3513 => x"5e",
  3514 => x"5b",
  3515 => x"5c",
  3516 => x"0e",
  3517 => x"71",
  3518 => x"4b",
  3519 => x"c0",
  3520 => x"4c",
  3521 => x"13",
  3522 => x"4a",
  3523 => x"72",
  3524 => x"9a",
  3525 => x"02",
  3526 => x"ce",
  3527 => x"87",
  3528 => x"72",
  3529 => x"49",
  3530 => x"ff",
  3531 => x"dd",
  3532 => x"87",
  3533 => x"c1",
  3534 => x"84",
  3535 => x"13",
  3536 => x"4a",
  3537 => x"72",
  3538 => x"9a",
  3539 => x"05",
  3540 => x"f2",
  3541 => x"87",
  3542 => x"74",
  3543 => x"48",
  3544 => x"c2",
  3545 => x"87",
  3546 => x"26",
  3547 => x"4d",
  3548 => x"26",
  3549 => x"4c",
  3550 => x"26",
  3551 => x"4b",
  3552 => x"26",
  3553 => x"4f",
  3554 => x"0e",
  3555 => x"5e",
  3556 => x"5b",
  3557 => x"5c",
  3558 => x"5d",
  3559 => x"0e",
  3560 => x"1e",
  3561 => x"d4",
  3562 => x"66",
  3563 => x"4b",
  3564 => x"c0",
  3565 => x"4c",
  3566 => x"b7",
  3567 => x"ab",
  3568 => x"06",
  3569 => x"c1",
  3570 => x"ca",
  3571 => x"87",
  3572 => x"11",
  3573 => x"4a",
  3574 => x"c8",
  3575 => x"32",
  3576 => x"c1",
  3577 => x"8b",
  3578 => x"c0",
  3579 => x"b7",
  3580 => x"ab",
  3581 => x"06",
  3582 => x"c7",
  3583 => x"87",
  3584 => x"11",
  3585 => x"48",
  3586 => x"c4",
  3587 => x"a6",
  3588 => x"58",
  3589 => x"c2",
  3590 => x"87",
  3591 => x"c0",
  3592 => x"7e",
  3593 => x"6e",
  3594 => x"b2",
  3595 => x"c8",
  3596 => x"32",
  3597 => x"c1",
  3598 => x"8b",
  3599 => x"c0",
  3600 => x"b7",
  3601 => x"ab",
  3602 => x"06",
  3603 => x"c4",
  3604 => x"87",
  3605 => x"11",
  3606 => x"4d",
  3607 => x"c2",
  3608 => x"87",
  3609 => x"c0",
  3610 => x"4d",
  3611 => x"75",
  3612 => x"b2",
  3613 => x"c8",
  3614 => x"32",
  3615 => x"c1",
  3616 => x"8b",
  3617 => x"c0",
  3618 => x"b7",
  3619 => x"ab",
  3620 => x"06",
  3621 => x"c7",
  3622 => x"87",
  3623 => x"11",
  3624 => x"48",
  3625 => x"c4",
  3626 => x"a6",
  3627 => x"58",
  3628 => x"c2",
  3629 => x"87",
  3630 => x"c0",
  3631 => x"7e",
  3632 => x"6e",
  3633 => x"b2",
  3634 => x"72",
  3635 => x"a4",
  3636 => x"4c",
  3637 => x"c1",
  3638 => x"8b",
  3639 => x"c0",
  3640 => x"b7",
  3641 => x"ab",
  3642 => x"01",
  3643 => x"fe",
  3644 => x"f6",
  3645 => x"87",
  3646 => x"74",
  3647 => x"48",
  3648 => x"26",
  3649 => x"26",
  3650 => x"4d",
  3651 => x"26",
  3652 => x"4c",
  3653 => x"26",
  3654 => x"4b",
  3655 => x"26",
  3656 => x"4f",
  3657 => x"0e",
  3658 => x"5e",
  3659 => x"5b",
  3660 => x"5c",
  3661 => x"5d",
  3662 => x"0e",
  3663 => x"71",
  3664 => x"4b",
  3665 => x"73",
  3666 => x"4c",
  3667 => x"d0",
  3668 => x"66",
  3669 => x"48",
  3670 => x"c2",
  3671 => x"28",
  3672 => x"d4",
  3673 => x"a6",
  3674 => x"58",
  3675 => x"d0",
  3676 => x"66",
  3677 => x"49",
  3678 => x"48",
  3679 => x"c1",
  3680 => x"88",
  3681 => x"d4",
  3682 => x"a6",
  3683 => x"58",
  3684 => x"71",
  3685 => x"99",
  3686 => x"02",
  3687 => x"c1",
  3688 => x"c4",
  3689 => x"87",
  3690 => x"24",
  3691 => x"4d",
  3692 => x"c0",
  3693 => x"4b",
  3694 => x"75",
  3695 => x"4a",
  3696 => x"dc",
  3697 => x"2a",
  3698 => x"c0",
  3699 => x"f0",
  3700 => x"82",
  3701 => x"c0",
  3702 => x"f9",
  3703 => x"aa",
  3704 => x"06",
  3705 => x"c2",
  3706 => x"87",
  3707 => x"c7",
  3708 => x"82",
  3709 => x"72",
  3710 => x"49",
  3711 => x"fc",
  3712 => x"e8",
  3713 => x"87",
  3714 => x"c4",
  3715 => x"35",
  3716 => x"c1",
  3717 => x"83",
  3718 => x"c8",
  3719 => x"b7",
  3720 => x"ab",
  3721 => x"04",
  3722 => x"e2",
  3723 => x"87",
  3724 => x"c0",
  3725 => x"e0",
  3726 => x"49",
  3727 => x"fc",
  3728 => x"d8",
  3729 => x"87",
  3730 => x"d0",
  3731 => x"66",
  3732 => x"49",
  3733 => x"c3",
  3734 => x"99",
  3735 => x"05",
  3736 => x"c5",
  3737 => x"87",
  3738 => x"ca",
  3739 => x"49",
  3740 => x"fc",
  3741 => x"cb",
  3742 => x"87",
  3743 => x"d0",
  3744 => x"66",
  3745 => x"49",
  3746 => x"48",
  3747 => x"c1",
  3748 => x"88",
  3749 => x"d4",
  3750 => x"a6",
  3751 => x"58",
  3752 => x"71",
  3753 => x"99",
  3754 => x"05",
  3755 => x"fe",
  3756 => x"fc",
  3757 => x"87",
  3758 => x"ca",
  3759 => x"49",
  3760 => x"fb",
  3761 => x"f7",
  3762 => x"87",
  3763 => x"26",
  3764 => x"4d",
  3765 => x"26",
  3766 => x"4c",
  3767 => x"26",
  3768 => x"4b",
  3769 => x"26",
  3770 => x"4f",
  3771 => x"0e",
  3772 => x"5e",
  3773 => x"5b",
  3774 => x"5c",
  3775 => x"5d",
  3776 => x"0e",
  3777 => x"fc",
  3778 => x"86",
  3779 => x"71",
  3780 => x"4a",
  3781 => x"c0",
  3782 => x"e0",
  3783 => x"66",
  3784 => x"4c",
  3785 => x"c1",
  3786 => x"d1",
  3787 => x"da",
  3788 => x"4b",
  3789 => x"c0",
  3790 => x"7e",
  3791 => x"72",
  3792 => x"9a",
  3793 => x"05",
  3794 => x"ce",
  3795 => x"87",
  3796 => x"c1",
  3797 => x"d1",
  3798 => x"db",
  3799 => x"4b",
  3800 => x"c1",
  3801 => x"d1",
  3802 => x"da",
  3803 => x"48",
  3804 => x"c0",
  3805 => x"f0",
  3806 => x"50",
  3807 => x"c1",
  3808 => x"d2",
  3809 => x"87",
  3810 => x"72",
  3811 => x"9a",
  3812 => x"02",
  3813 => x"c0",
  3814 => x"e9",
  3815 => x"87",
  3816 => x"d4",
  3817 => x"66",
  3818 => x"4d",
  3819 => x"72",
  3820 => x"1e",
  3821 => x"72",
  3822 => x"49",
  3823 => x"75",
  3824 => x"4a",
  3825 => x"ca",
  3826 => x"cf",
  3827 => x"87",
  3828 => x"26",
  3829 => x"4a",
  3830 => x"c0",
  3831 => x"fd",
  3832 => x"e5",
  3833 => x"81",
  3834 => x"11",
  3835 => x"53",
  3836 => x"71",
  3837 => x"1e",
  3838 => x"72",
  3839 => x"49",
  3840 => x"75",
  3841 => x"4a",
  3842 => x"c9",
  3843 => x"fe",
  3844 => x"87",
  3845 => x"70",
  3846 => x"4a",
  3847 => x"26",
  3848 => x"49",
  3849 => x"c1",
  3850 => x"8c",
  3851 => x"72",
  3852 => x"9a",
  3853 => x"05",
  3854 => x"ff",
  3855 => x"da",
  3856 => x"87",
  3857 => x"c0",
  3858 => x"b7",
  3859 => x"ac",
  3860 => x"06",
  3861 => x"dd",
  3862 => x"87",
  3863 => x"c0",
  3864 => x"e4",
  3865 => x"66",
  3866 => x"02",
  3867 => x"c5",
  3868 => x"87",
  3869 => x"c0",
  3870 => x"f0",
  3871 => x"4a",
  3872 => x"c3",
  3873 => x"87",
  3874 => x"c0",
  3875 => x"e0",
  3876 => x"4a",
  3877 => x"73",
  3878 => x"0a",
  3879 => x"97",
  3880 => x"7a",
  3881 => x"0a",
  3882 => x"c1",
  3883 => x"83",
  3884 => x"8c",
  3885 => x"c0",
  3886 => x"b7",
  3887 => x"ac",
  3888 => x"01",
  3889 => x"ff",
  3890 => x"e3",
  3891 => x"87",
  3892 => x"c1",
  3893 => x"d1",
  3894 => x"da",
  3895 => x"ab",
  3896 => x"02",
  3897 => x"de",
  3898 => x"87",
  3899 => x"d8",
  3900 => x"66",
  3901 => x"4c",
  3902 => x"dc",
  3903 => x"66",
  3904 => x"1e",
  3905 => x"c1",
  3906 => x"8b",
  3907 => x"97",
  3908 => x"6b",
  3909 => x"49",
  3910 => x"74",
  3911 => x"0f",
  3912 => x"c4",
  3913 => x"86",
  3914 => x"6e",
  3915 => x"48",
  3916 => x"c1",
  3917 => x"80",
  3918 => x"c4",
  3919 => x"a6",
  3920 => x"58",
  3921 => x"c1",
  3922 => x"d1",
  3923 => x"da",
  3924 => x"ab",
  3925 => x"05",
  3926 => x"ff",
  3927 => x"e5",
  3928 => x"87",
  3929 => x"6e",
  3930 => x"48",
  3931 => x"fc",
  3932 => x"8e",
  3933 => x"26",
  3934 => x"4d",
  3935 => x"26",
  3936 => x"4c",
  3937 => x"26",
  3938 => x"4b",
  3939 => x"26",
  3940 => x"4f",
  3941 => x"30",
  3942 => x"31",
  3943 => x"32",
  3944 => x"33",
  3945 => x"34",
  3946 => x"35",
  3947 => x"36",
  3948 => x"37",
  3949 => x"38",
  3950 => x"39",
  3951 => x"41",
  3952 => x"42",
  3953 => x"43",
  3954 => x"44",
  3955 => x"45",
  3956 => x"46",
  3957 => x"00",
  3958 => x"0e",
  3959 => x"5e",
  3960 => x"5b",
  3961 => x"5c",
  3962 => x"5d",
  3963 => x"0e",
  3964 => x"71",
  3965 => x"4b",
  3966 => x"ff",
  3967 => x"4d",
  3968 => x"13",
  3969 => x"4c",
  3970 => x"74",
  3971 => x"9c",
  3972 => x"02",
  3973 => x"d8",
  3974 => x"87",
  3975 => x"c1",
  3976 => x"85",
  3977 => x"d4",
  3978 => x"66",
  3979 => x"1e",
  3980 => x"74",
  3981 => x"49",
  3982 => x"d4",
  3983 => x"66",
  3984 => x"0f",
  3985 => x"c4",
  3986 => x"86",
  3987 => x"74",
  3988 => x"a8",
  3989 => x"05",
  3990 => x"c7",
  3991 => x"87",
  3992 => x"13",
  3993 => x"4c",
  3994 => x"74",
  3995 => x"9c",
  3996 => x"05",
  3997 => x"e8",
  3998 => x"87",
  3999 => x"75",
  4000 => x"48",
  4001 => x"26",
  4002 => x"4d",
  4003 => x"26",
  4004 => x"4c",
  4005 => x"26",
  4006 => x"4b",
  4007 => x"26",
  4008 => x"4f",
  4009 => x"0e",
  4010 => x"5e",
  4011 => x"5b",
  4012 => x"5c",
  4013 => x"5d",
  4014 => x"0e",
  4015 => x"e8",
  4016 => x"86",
  4017 => x"c4",
  4018 => x"a6",
  4019 => x"59",
  4020 => x"c0",
  4021 => x"e8",
  4022 => x"66",
  4023 => x"4d",
  4024 => x"c0",
  4025 => x"4c",
  4026 => x"c8",
  4027 => x"a6",
  4028 => x"48",
  4029 => x"c0",
  4030 => x"78",
  4031 => x"6e",
  4032 => x"97",
  4033 => x"bf",
  4034 => x"4b",
  4035 => x"6e",
  4036 => x"48",
  4037 => x"c1",
  4038 => x"80",
  4039 => x"c4",
  4040 => x"a6",
  4041 => x"58",
  4042 => x"73",
  4043 => x"9b",
  4044 => x"02",
  4045 => x"c6",
  4046 => x"d3",
  4047 => x"87",
  4048 => x"c8",
  4049 => x"66",
  4050 => x"02",
  4051 => x"c5",
  4052 => x"db",
  4053 => x"87",
  4054 => x"cc",
  4055 => x"a6",
  4056 => x"48",
  4057 => x"c0",
  4058 => x"78",
  4059 => x"fc",
  4060 => x"80",
  4061 => x"c0",
  4062 => x"78",
  4063 => x"73",
  4064 => x"4a",
  4065 => x"c0",
  4066 => x"e0",
  4067 => x"8a",
  4068 => x"02",
  4069 => x"c3",
  4070 => x"c6",
  4071 => x"87",
  4072 => x"c3",
  4073 => x"8a",
  4074 => x"02",
  4075 => x"c3",
  4076 => x"c0",
  4077 => x"87",
  4078 => x"c2",
  4079 => x"8a",
  4080 => x"02",
  4081 => x"c2",
  4082 => x"e8",
  4083 => x"87",
  4084 => x"c2",
  4085 => x"8a",
  4086 => x"02",
  4087 => x"c2",
  4088 => x"f4",
  4089 => x"87",
  4090 => x"c4",
  4091 => x"8a",
  4092 => x"02",
  4093 => x"c2",
  4094 => x"ee",
  4095 => x"87",
  4096 => x"c2",
  4097 => x"8a",
  4098 => x"02",
  4099 => x"c2",
  4100 => x"e8",
  4101 => x"87",
  4102 => x"c3",
  4103 => x"8a",
  4104 => x"02",
  4105 => x"c2",
  4106 => x"ea",
  4107 => x"87",
  4108 => x"d4",
  4109 => x"8a",
  4110 => x"02",
  4111 => x"c0",
  4112 => x"f6",
  4113 => x"87",
  4114 => x"d4",
  4115 => x"8a",
  4116 => x"02",
  4117 => x"c1",
  4118 => x"c0",
  4119 => x"87",
  4120 => x"ca",
  4121 => x"8a",
  4122 => x"02",
  4123 => x"c0",
  4124 => x"f2",
  4125 => x"87",
  4126 => x"c1",
  4127 => x"8a",
  4128 => x"02",
  4129 => x"c1",
  4130 => x"e1",
  4131 => x"87",
  4132 => x"c1",
  4133 => x"8a",
  4134 => x"02",
  4135 => x"df",
  4136 => x"87",
  4137 => x"c8",
  4138 => x"8a",
  4139 => x"02",
  4140 => x"c1",
  4141 => x"ce",
  4142 => x"87",
  4143 => x"c4",
  4144 => x"8a",
  4145 => x"02",
  4146 => x"c0",
  4147 => x"e3",
  4148 => x"87",
  4149 => x"c3",
  4150 => x"8a",
  4151 => x"02",
  4152 => x"c0",
  4153 => x"e5",
  4154 => x"87",
  4155 => x"c2",
  4156 => x"8a",
  4157 => x"02",
  4158 => x"c8",
  4159 => x"87",
  4160 => x"c3",
  4161 => x"8a",
  4162 => x"02",
  4163 => x"d3",
  4164 => x"87",
  4165 => x"c1",
  4166 => x"fa",
  4167 => x"87",
  4168 => x"cc",
  4169 => x"a6",
  4170 => x"48",
  4171 => x"ca",
  4172 => x"78",
  4173 => x"c2",
  4174 => x"d2",
  4175 => x"87",
  4176 => x"cc",
  4177 => x"a6",
  4178 => x"48",
  4179 => x"c2",
  4180 => x"78",
  4181 => x"c2",
  4182 => x"ca",
  4183 => x"87",
  4184 => x"cc",
  4185 => x"a6",
  4186 => x"48",
  4187 => x"d0",
  4188 => x"78",
  4189 => x"c2",
  4190 => x"c2",
  4191 => x"87",
  4192 => x"c0",
  4193 => x"f0",
  4194 => x"66",
  4195 => x"1e",
  4196 => x"c0",
  4197 => x"f0",
  4198 => x"66",
  4199 => x"1e",
  4200 => x"c4",
  4201 => x"85",
  4202 => x"75",
  4203 => x"4a",
  4204 => x"c4",
  4205 => x"8a",
  4206 => x"6a",
  4207 => x"49",
  4208 => x"fc",
  4209 => x"c3",
  4210 => x"87",
  4211 => x"c8",
  4212 => x"86",
  4213 => x"70",
  4214 => x"49",
  4215 => x"71",
  4216 => x"a4",
  4217 => x"4c",
  4218 => x"c1",
  4219 => x"e5",
  4220 => x"87",
  4221 => x"c8",
  4222 => x"a6",
  4223 => x"48",
  4224 => x"c1",
  4225 => x"78",
  4226 => x"c1",
  4227 => x"dd",
  4228 => x"87",
  4229 => x"c0",
  4230 => x"f0",
  4231 => x"66",
  4232 => x"1e",
  4233 => x"c4",
  4234 => x"85",
  4235 => x"75",
  4236 => x"4a",
  4237 => x"c4",
  4238 => x"8a",
  4239 => x"6a",
  4240 => x"49",
  4241 => x"c0",
  4242 => x"f0",
  4243 => x"66",
  4244 => x"0f",
  4245 => x"c4",
  4246 => x"86",
  4247 => x"c1",
  4248 => x"84",
  4249 => x"c1",
  4250 => x"c6",
  4251 => x"87",
  4252 => x"c0",
  4253 => x"f0",
  4254 => x"66",
  4255 => x"1e",
  4256 => x"c0",
  4257 => x"e5",
  4258 => x"49",
  4259 => x"c0",
  4260 => x"f0",
  4261 => x"66",
  4262 => x"0f",
  4263 => x"c4",
  4264 => x"86",
  4265 => x"c1",
  4266 => x"84",
  4267 => x"c0",
  4268 => x"f4",
  4269 => x"87",
  4270 => x"c8",
  4271 => x"a6",
  4272 => x"48",
  4273 => x"c1",
  4274 => x"78",
  4275 => x"c0",
  4276 => x"ec",
  4277 => x"87",
  4278 => x"d0",
  4279 => x"a6",
  4280 => x"48",
  4281 => x"c1",
  4282 => x"78",
  4283 => x"f8",
  4284 => x"80",
  4285 => x"c1",
  4286 => x"78",
  4287 => x"c0",
  4288 => x"e0",
  4289 => x"87",
  4290 => x"c0",
  4291 => x"f0",
  4292 => x"ab",
  4293 => x"06",
  4294 => x"da",
  4295 => x"87",
  4296 => x"c0",
  4297 => x"f9",
  4298 => x"ab",
  4299 => x"03",
  4300 => x"d4",
  4301 => x"87",
  4302 => x"d4",
  4303 => x"66",
  4304 => x"49",
  4305 => x"ca",
  4306 => x"91",
  4307 => x"73",
  4308 => x"4a",
  4309 => x"c0",
  4310 => x"f0",
  4311 => x"8a",
  4312 => x"d4",
  4313 => x"a6",
  4314 => x"48",
  4315 => x"72",
  4316 => x"a1",
  4317 => x"78",
  4318 => x"f4",
  4319 => x"80",
  4320 => x"c1",
  4321 => x"78",
  4322 => x"cc",
  4323 => x"66",
  4324 => x"02",
  4325 => x"c1",
  4326 => x"ea",
  4327 => x"87",
  4328 => x"c4",
  4329 => x"85",
  4330 => x"75",
  4331 => x"49",
  4332 => x"c4",
  4333 => x"89",
  4334 => x"a6",
  4335 => x"48",
  4336 => x"69",
  4337 => x"78",
  4338 => x"c1",
  4339 => x"e4",
  4340 => x"ab",
  4341 => x"05",
  4342 => x"d8",
  4343 => x"87",
  4344 => x"c4",
  4345 => x"66",
  4346 => x"48",
  4347 => x"c0",
  4348 => x"b7",
  4349 => x"a8",
  4350 => x"03",
  4351 => x"cf",
  4352 => x"87",
  4353 => x"c0",
  4354 => x"ed",
  4355 => x"49",
  4356 => x"f2",
  4357 => x"e3",
  4358 => x"87",
  4359 => x"c4",
  4360 => x"66",
  4361 => x"48",
  4362 => x"c0",
  4363 => x"08",
  4364 => x"88",
  4365 => x"c8",
  4366 => x"a6",
  4367 => x"58",
  4368 => x"d0",
  4369 => x"66",
  4370 => x"1e",
  4371 => x"d8",
  4372 => x"66",
  4373 => x"1e",
  4374 => x"c0",
  4375 => x"f8",
  4376 => x"66",
  4377 => x"1e",
  4378 => x"c0",
  4379 => x"f8",
  4380 => x"66",
  4381 => x"1e",
  4382 => x"dc",
  4383 => x"66",
  4384 => x"1e",
  4385 => x"d8",
  4386 => x"66",
  4387 => x"49",
  4388 => x"f6",
  4389 => x"d4",
  4390 => x"87",
  4391 => x"d4",
  4392 => x"86",
  4393 => x"70",
  4394 => x"49",
  4395 => x"71",
  4396 => x"a4",
  4397 => x"4c",
  4398 => x"c0",
  4399 => x"e1",
  4400 => x"87",
  4401 => x"c0",
  4402 => x"e5",
  4403 => x"ab",
  4404 => x"05",
  4405 => x"cf",
  4406 => x"87",
  4407 => x"d0",
  4408 => x"a6",
  4409 => x"48",
  4410 => x"c0",
  4411 => x"78",
  4412 => x"c4",
  4413 => x"80",
  4414 => x"c0",
  4415 => x"78",
  4416 => x"f4",
  4417 => x"80",
  4418 => x"c1",
  4419 => x"78",
  4420 => x"cc",
  4421 => x"87",
  4422 => x"c0",
  4423 => x"f0",
  4424 => x"66",
  4425 => x"1e",
  4426 => x"73",
  4427 => x"49",
  4428 => x"c0",
  4429 => x"f0",
  4430 => x"66",
  4431 => x"0f",
  4432 => x"c4",
  4433 => x"86",
  4434 => x"6e",
  4435 => x"97",
  4436 => x"bf",
  4437 => x"4b",
  4438 => x"6e",
  4439 => x"48",
  4440 => x"c1",
  4441 => x"80",
  4442 => x"c4",
  4443 => x"a6",
  4444 => x"58",
  4445 => x"73",
  4446 => x"9b",
  4447 => x"05",
  4448 => x"f9",
  4449 => x"ed",
  4450 => x"87",
  4451 => x"74",
  4452 => x"48",
  4453 => x"e8",
  4454 => x"8e",
  4455 => x"26",
  4456 => x"4d",
  4457 => x"26",
  4458 => x"4c",
  4459 => x"26",
  4460 => x"4b",
  4461 => x"26",
  4462 => x"4f",
  4463 => x"1e",
  4464 => x"c0",
  4465 => x"1e",
  4466 => x"c0",
  4467 => x"f6",
  4468 => x"ea",
  4469 => x"1e",
  4470 => x"d0",
  4471 => x"a6",
  4472 => x"1e",
  4473 => x"d0",
  4474 => x"66",
  4475 => x"49",
  4476 => x"f8",
  4477 => x"ea",
  4478 => x"87",
  4479 => x"f4",
  4480 => x"8e",
  4481 => x"26",
  4482 => x"4f",
  4483 => x"1e",
  4484 => x"73",
  4485 => x"1e",
  4486 => x"72",
  4487 => x"9a",
  4488 => x"02",
  4489 => x"c0",
  4490 => x"e7",
  4491 => x"87",
  4492 => x"c0",
  4493 => x"48",
  4494 => x"c1",
  4495 => x"4b",
  4496 => x"72",
  4497 => x"a9",
  4498 => x"06",
  4499 => x"d1",
  4500 => x"87",
  4501 => x"72",
  4502 => x"82",
  4503 => x"06",
  4504 => x"c9",
  4505 => x"87",
  4506 => x"73",
  4507 => x"83",
  4508 => x"72",
  4509 => x"a9",
  4510 => x"01",
  4511 => x"f4",
  4512 => x"87",
  4513 => x"c3",
  4514 => x"87",
  4515 => x"c1",
  4516 => x"b2",
  4517 => x"3a",
  4518 => x"72",
  4519 => x"a9",
  4520 => x"03",
  4521 => x"89",
  4522 => x"73",
  4523 => x"80",
  4524 => x"07",
  4525 => x"c1",
  4526 => x"2a",
  4527 => x"2b",
  4528 => x"05",
  4529 => x"f3",
  4530 => x"87",
  4531 => x"26",
  4532 => x"4b",
  4533 => x"26",
  4534 => x"4f",
  4535 => x"1e",
  4536 => x"75",
  4537 => x"1e",
  4538 => x"c4",
  4539 => x"4d",
  4540 => x"71",
  4541 => x"b7",
  4542 => x"a1",
  4543 => x"04",
  4544 => x"ff",
  4545 => x"b9",
  4546 => x"c1",
  4547 => x"81",
  4548 => x"c3",
  4549 => x"bd",
  4550 => x"07",
  4551 => x"72",
  4552 => x"b7",
  4553 => x"a2",
  4554 => x"04",
  4555 => x"ff",
  4556 => x"ba",
  4557 => x"c1",
  4558 => x"82",
  4559 => x"c1",
  4560 => x"bd",
  4561 => x"07",
  4562 => x"fe",
  4563 => x"ee",
  4564 => x"87",
  4565 => x"c1",
  4566 => x"2d",
  4567 => x"04",
  4568 => x"ff",
  4569 => x"b8",
  4570 => x"c1",
  4571 => x"80",
  4572 => x"07",
  4573 => x"2d",
  4574 => x"04",
  4575 => x"ff",
  4576 => x"b9",
  4577 => x"c1",
  4578 => x"81",
  4579 => x"07",
  4580 => x"26",
  4581 => x"4d",
  4582 => x"26",
  4583 => x"4f",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;

