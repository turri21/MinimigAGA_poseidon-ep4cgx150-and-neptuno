library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"01",
     1 => x"da",
     2 => x"87",
     3 => x"04",
     4 => x"dd",
     5 => x"87",
     6 => x"0e",
     7 => x"58",
     8 => x"5e",
     9 => x"59",
    10 => x"5a",
    11 => x"0e",
    12 => x"27",
    13 => x"00",
    14 => x"00",
    15 => x"00",
    16 => x"2c",
    17 => x"0f",
    18 => x"26",
    19 => x"4a",
    20 => x"26",
    21 => x"49",
    22 => x"26",
    23 => x"48",
    24 => x"ff",
    25 => x"80",
    26 => x"26",
    27 => x"08",
    28 => x"4f",
    29 => x"27",
    30 => x"00",
    31 => x"00",
    32 => x"00",
    33 => x"2d",
    34 => x"4f",
    35 => x"27",
    36 => x"00",
    37 => x"00",
    38 => x"00",
    39 => x"29",
    40 => x"4f",
    41 => x"00",
    42 => x"fd",
    43 => x"87",
    44 => x"4f",
    45 => x"c1",
    46 => x"cb",
    47 => x"fc",
    48 => x"4e",
    49 => x"c9",
    50 => x"c0",
    51 => x"86",
    52 => x"c1",
    53 => x"cb",
    54 => x"fc",
    55 => x"49",
    56 => x"c1",
    57 => x"c2",
    58 => x"d8",
    59 => x"48",
    60 => x"89",
    61 => x"d0",
    62 => x"89",
    63 => x"03",
    64 => x"c0",
    65 => x"40",
    66 => x"40",
    67 => x"40",
    68 => x"40",
    69 => x"f6",
    70 => x"87",
    71 => x"d0",
    72 => x"81",
    73 => x"05",
    74 => x"c0",
    75 => x"50",
    76 => x"c1",
    77 => x"89",
    78 => x"05",
    79 => x"f9",
    80 => x"87",
    81 => x"c1",
    82 => x"c2",
    83 => x"d7",
    84 => x"4d",
    85 => x"c1",
    86 => x"c2",
    87 => x"d7",
    88 => x"4c",
    89 => x"74",
    90 => x"ad",
    91 => x"02",
    92 => x"c4",
    93 => x"87",
    94 => x"24",
    95 => x"0f",
    96 => x"f7",
    97 => x"87",
    98 => x"c1",
    99 => x"c0",
   100 => x"87",
   101 => x"c1",
   102 => x"c2",
   103 => x"d7",
   104 => x"4d",
   105 => x"c1",
   106 => x"c2",
   107 => x"d7",
   108 => x"4c",
   109 => x"74",
   110 => x"ad",
   111 => x"02",
   112 => x"c6",
   113 => x"87",
   114 => x"c4",
   115 => x"8c",
   116 => x"6c",
   117 => x"0f",
   118 => x"f5",
   119 => x"87",
   120 => x"00",
   121 => x"fd",
   122 => x"87",
   123 => x"1e",
   124 => x"73",
   125 => x"1e",
   126 => x"c2",
   127 => x"c0",
   128 => x"c0",
   129 => x"4b",
   130 => x"73",
   131 => x"0f",
   132 => x"c4",
   133 => x"87",
   134 => x"26",
   135 => x"4d",
   136 => x"26",
   137 => x"4c",
   138 => x"26",
   139 => x"4b",
   140 => x"26",
   141 => x"4f",
   142 => x"1e",
   143 => x"e5",
   144 => x"48",
   145 => x"c0",
   146 => x"e0",
   147 => x"50",
   148 => x"e5",
   149 => x"48",
   150 => x"c0",
   151 => x"e1",
   152 => x"50",
   153 => x"e5",
   154 => x"48",
   155 => x"c0",
   156 => x"e0",
   157 => x"50",
   158 => x"e5",
   159 => x"48",
   160 => x"c0",
   161 => x"e1",
   162 => x"50",
   163 => x"26",
   164 => x"4f",
   165 => x"1e",
   166 => x"73",
   167 => x"1e",
   168 => x"c4",
   169 => x"fa",
   170 => x"49",
   171 => x"c0",
   172 => x"f0",
   173 => x"e0",
   174 => x"87",
   175 => x"c0",
   176 => x"fc",
   177 => x"c0",
   178 => x"4b",
   179 => x"cf",
   180 => x"da",
   181 => x"87",
   182 => x"70",
   183 => x"98",
   184 => x"02",
   185 => x"c0",
   186 => x"f4",
   187 => x"87",
   188 => x"c0",
   189 => x"ff",
   190 => x"f0",
   191 => x"4b",
   192 => x"c4",
   193 => x"e3",
   194 => x"49",
   195 => x"c0",
   196 => x"f0",
   197 => x"c8",
   198 => x"87",
   199 => x"d5",
   200 => x"cd",
   201 => x"87",
   202 => x"70",
   203 => x"98",
   204 => x"02",
   205 => x"da",
   206 => x"87",
   207 => x"c3",
   208 => x"f0",
   209 => x"4b",
   210 => x"c2",
   211 => x"c0",
   212 => x"c0",
   213 => x"1e",
   214 => x"c3",
   215 => x"fb",
   216 => x"49",
   217 => x"c0",
   218 => x"ec",
   219 => x"ff",
   220 => x"87",
   221 => x"c4",
   222 => x"86",
   223 => x"70",
   224 => x"98",
   225 => x"02",
   226 => x"cc",
   227 => x"87",
   228 => x"fe",
   229 => x"d4",
   230 => x"87",
   231 => x"c7",
   232 => x"87",
   233 => x"c4",
   234 => x"c7",
   235 => x"49",
   236 => x"c0",
   237 => x"ef",
   238 => x"df",
   239 => x"87",
   240 => x"73",
   241 => x"49",
   242 => x"fe",
   243 => x"d9",
   244 => x"87",
   245 => x"fe",
   246 => x"f0",
   247 => x"87",
   248 => x"fe",
   249 => x"cf",
   250 => x"87",
   251 => x"38",
   252 => x"33",
   253 => x"32",
   254 => x"4f",
   255 => x"53",
   256 => x"44",
   257 => x"41",
   258 => x"42",
   259 => x"42",
   260 => x"49",
   261 => x"4e",
   262 => x"00",
   263 => x"55",
   264 => x"6e",
   265 => x"61",
   266 => x"62",
   267 => x"6c",
   268 => x"65",
   269 => x"20",
   270 => x"74",
   271 => x"6f",
   272 => x"20",
   273 => x"6c",
   274 => x"6f",
   275 => x"63",
   276 => x"61",
   277 => x"74",
   278 => x"65",
   279 => x"20",
   280 => x"70",
   281 => x"61",
   282 => x"72",
   283 => x"74",
   284 => x"69",
   285 => x"74",
   286 => x"69",
   287 => x"6f",
   288 => x"6e",
   289 => x"0a",
   290 => x"00",
   291 => x"48",
   292 => x"75",
   293 => x"6e",
   294 => x"74",
   295 => x"69",
   296 => x"6e",
   297 => x"67",
   298 => x"20",
   299 => x"66",
   300 => x"6f",
   301 => x"72",
   302 => x"20",
   303 => x"70",
   304 => x"61",
   305 => x"72",
   306 => x"74",
   307 => x"69",
   308 => x"74",
   309 => x"69",
   310 => x"6f",
   311 => x"6e",
   312 => x"0a",
   313 => x"00",
   314 => x"49",
   315 => x"6e",
   316 => x"69",
   317 => x"74",
   318 => x"69",
   319 => x"61",
   320 => x"6c",
   321 => x"69",
   322 => x"7a",
   323 => x"69",
   324 => x"6e",
   325 => x"67",
   326 => x"20",
   327 => x"53",
   328 => x"44",
   329 => x"20",
   330 => x"63",
   331 => x"61",
   332 => x"72",
   333 => x"64",
   334 => x"0a",
   335 => x"00",
   336 => x"1e",
   337 => x"e4",
   338 => x"86",
   339 => x"e1",
   340 => x"48",
   341 => x"c3",
   342 => x"ff",
   343 => x"50",
   344 => x"e1",
   345 => x"97",
   346 => x"bf",
   347 => x"48",
   348 => x"c4",
   349 => x"a6",
   350 => x"58",
   351 => x"6e",
   352 => x"49",
   353 => x"c3",
   354 => x"ff",
   355 => x"99",
   356 => x"e1",
   357 => x"48",
   358 => x"c3",
   359 => x"ff",
   360 => x"50",
   361 => x"c8",
   362 => x"31",
   363 => x"e1",
   364 => x"97",
   365 => x"bf",
   366 => x"48",
   367 => x"c8",
   368 => x"a6",
   369 => x"58",
   370 => x"c4",
   371 => x"66",
   372 => x"48",
   373 => x"c3",
   374 => x"ff",
   375 => x"98",
   376 => x"cc",
   377 => x"a6",
   378 => x"58",
   379 => x"c8",
   380 => x"66",
   381 => x"b1",
   382 => x"e1",
   383 => x"48",
   384 => x"c3",
   385 => x"ff",
   386 => x"50",
   387 => x"c8",
   388 => x"31",
   389 => x"e1",
   390 => x"97",
   391 => x"bf",
   392 => x"48",
   393 => x"d0",
   394 => x"a6",
   395 => x"58",
   396 => x"cc",
   397 => x"66",
   398 => x"48",
   399 => x"c3",
   400 => x"ff",
   401 => x"98",
   402 => x"d4",
   403 => x"a6",
   404 => x"58",
   405 => x"d0",
   406 => x"66",
   407 => x"b1",
   408 => x"e1",
   409 => x"48",
   410 => x"c3",
   411 => x"ff",
   412 => x"50",
   413 => x"c8",
   414 => x"31",
   415 => x"e1",
   416 => x"97",
   417 => x"bf",
   418 => x"48",
   419 => x"d8",
   420 => x"a6",
   421 => x"58",
   422 => x"d4",
   423 => x"66",
   424 => x"48",
   425 => x"c3",
   426 => x"ff",
   427 => x"98",
   428 => x"dc",
   429 => x"a6",
   430 => x"58",
   431 => x"d8",
   432 => x"66",
   433 => x"b1",
   434 => x"71",
   435 => x"48",
   436 => x"e4",
   437 => x"8e",
   438 => x"26",
   439 => x"4f",
   440 => x"0e",
   441 => x"5e",
   442 => x"5b",
   443 => x"5c",
   444 => x"0e",
   445 => x"1e",
   446 => x"71",
   447 => x"4a",
   448 => x"72",
   449 => x"49",
   450 => x"c3",
   451 => x"ff",
   452 => x"99",
   453 => x"e1",
   454 => x"09",
   455 => x"97",
   456 => x"79",
   457 => x"09",
   458 => x"c1",
   459 => x"c2",
   460 => x"d8",
   461 => x"bf",
   462 => x"05",
   463 => x"c8",
   464 => x"87",
   465 => x"d0",
   466 => x"66",
   467 => x"48",
   468 => x"c9",
   469 => x"30",
   470 => x"d4",
   471 => x"a6",
   472 => x"58",
   473 => x"d0",
   474 => x"66",
   475 => x"49",
   476 => x"d8",
   477 => x"29",
   478 => x"c3",
   479 => x"ff",
   480 => x"99",
   481 => x"e1",
   482 => x"09",
   483 => x"97",
   484 => x"79",
   485 => x"09",
   486 => x"d0",
   487 => x"66",
   488 => x"49",
   489 => x"d0",
   490 => x"29",
   491 => x"c3",
   492 => x"ff",
   493 => x"99",
   494 => x"e1",
   495 => x"09",
   496 => x"97",
   497 => x"79",
   498 => x"09",
   499 => x"d0",
   500 => x"66",
   501 => x"49",
   502 => x"c8",
   503 => x"29",
   504 => x"c3",
   505 => x"ff",
   506 => x"99",
   507 => x"e1",
   508 => x"09",
   509 => x"97",
   510 => x"79",
   511 => x"09",
   512 => x"d0",
   513 => x"66",
   514 => x"49",
   515 => x"c3",
   516 => x"ff",
   517 => x"99",
   518 => x"e1",
   519 => x"09",
   520 => x"97",
   521 => x"79",
   522 => x"09",
   523 => x"72",
   524 => x"49",
   525 => x"d0",
   526 => x"29",
   527 => x"c3",
   528 => x"ff",
   529 => x"99",
   530 => x"e1",
   531 => x"09",
   532 => x"97",
   533 => x"79",
   534 => x"09",
   535 => x"97",
   536 => x"bf",
   537 => x"48",
   538 => x"c4",
   539 => x"a6",
   540 => x"58",
   541 => x"6e",
   542 => x"4b",
   543 => x"c3",
   544 => x"ff",
   545 => x"9b",
   546 => x"c9",
   547 => x"f0",
   548 => x"ff",
   549 => x"4c",
   550 => x"c3",
   551 => x"ff",
   552 => x"ab",
   553 => x"05",
   554 => x"dc",
   555 => x"87",
   556 => x"e1",
   557 => x"48",
   558 => x"c3",
   559 => x"ff",
   560 => x"50",
   561 => x"e1",
   562 => x"97",
   563 => x"bf",
   564 => x"48",
   565 => x"c4",
   566 => x"a6",
   567 => x"58",
   568 => x"6e",
   569 => x"4b",
   570 => x"c3",
   571 => x"ff",
   572 => x"9b",
   573 => x"c1",
   574 => x"8c",
   575 => x"02",
   576 => x"c6",
   577 => x"87",
   578 => x"c3",
   579 => x"ff",
   580 => x"ab",
   581 => x"02",
   582 => x"e4",
   583 => x"87",
   584 => x"73",
   585 => x"4a",
   586 => x"c4",
   587 => x"b7",
   588 => x"2a",
   589 => x"c0",
   590 => x"f0",
   591 => x"a2",
   592 => x"49",
   593 => x"c0",
   594 => x"e9",
   595 => x"f0",
   596 => x"87",
   597 => x"73",
   598 => x"4a",
   599 => x"cf",
   600 => x"9a",
   601 => x"c0",
   602 => x"f0",
   603 => x"a2",
   604 => x"49",
   605 => x"c0",
   606 => x"e9",
   607 => x"e4",
   608 => x"87",
   609 => x"73",
   610 => x"48",
   611 => x"26",
   612 => x"c2",
   613 => x"87",
   614 => x"26",
   615 => x"4d",
   616 => x"26",
   617 => x"4c",
   618 => x"26",
   619 => x"4b",
   620 => x"26",
   621 => x"4f",
   622 => x"1e",
   623 => x"c0",
   624 => x"49",
   625 => x"e1",
   626 => x"48",
   627 => x"c3",
   628 => x"ff",
   629 => x"50",
   630 => x"c1",
   631 => x"81",
   632 => x"c3",
   633 => x"c8",
   634 => x"b7",
   635 => x"a9",
   636 => x"04",
   637 => x"f2",
   638 => x"87",
   639 => x"26",
   640 => x"4f",
   641 => x"1e",
   642 => x"73",
   643 => x"1e",
   644 => x"e8",
   645 => x"87",
   646 => x"c4",
   647 => x"f8",
   648 => x"df",
   649 => x"4b",
   650 => x"c0",
   651 => x"1e",
   652 => x"c0",
   653 => x"ff",
   654 => x"f0",
   655 => x"c1",
   656 => x"f7",
   657 => x"49",
   658 => x"fc",
   659 => x"e3",
   660 => x"87",
   661 => x"c4",
   662 => x"86",
   663 => x"c1",
   664 => x"a8",
   665 => x"05",
   666 => x"c0",
   667 => x"e8",
   668 => x"87",
   669 => x"e1",
   670 => x"48",
   671 => x"c3",
   672 => x"ff",
   673 => x"50",
   674 => x"c1",
   675 => x"c0",
   676 => x"c0",
   677 => x"c0",
   678 => x"c0",
   679 => x"c0",
   680 => x"1e",
   681 => x"c0",
   682 => x"e1",
   683 => x"f0",
   684 => x"c1",
   685 => x"e9",
   686 => x"49",
   687 => x"fc",
   688 => x"c6",
   689 => x"87",
   690 => x"c4",
   691 => x"86",
   692 => x"70",
   693 => x"98",
   694 => x"05",
   695 => x"c9",
   696 => x"87",
   697 => x"e1",
   698 => x"48",
   699 => x"c3",
   700 => x"ff",
   701 => x"50",
   702 => x"c1",
   703 => x"48",
   704 => x"cb",
   705 => x"87",
   706 => x"fe",
   707 => x"e9",
   708 => x"87",
   709 => x"c1",
   710 => x"8b",
   711 => x"05",
   712 => x"fe",
   713 => x"ff",
   714 => x"87",
   715 => x"c0",
   716 => x"48",
   717 => x"fe",
   718 => x"da",
   719 => x"87",
   720 => x"43",
   721 => x"4d",
   722 => x"44",
   723 => x"34",
   724 => x"31",
   725 => x"20",
   726 => x"25",
   727 => x"64",
   728 => x"0a",
   729 => x"00",
   730 => x"43",
   731 => x"4d",
   732 => x"44",
   733 => x"35",
   734 => x"35",
   735 => x"20",
   736 => x"25",
   737 => x"64",
   738 => x"0a",
   739 => x"00",
   740 => x"43",
   741 => x"4d",
   742 => x"44",
   743 => x"34",
   744 => x"31",
   745 => x"20",
   746 => x"25",
   747 => x"64",
   748 => x"0a",
   749 => x"00",
   750 => x"43",
   751 => x"4d",
   752 => x"44",
   753 => x"35",
   754 => x"35",
   755 => x"20",
   756 => x"25",
   757 => x"64",
   758 => x"0a",
   759 => x"00",
   760 => x"69",
   761 => x"6e",
   762 => x"69",
   763 => x"74",
   764 => x"20",
   765 => x"25",
   766 => x"64",
   767 => x"0a",
   768 => x"20",
   769 => x"20",
   770 => x"00",
   771 => x"69",
   772 => x"6e",
   773 => x"69",
   774 => x"74",
   775 => x"20",
   776 => x"25",
   777 => x"64",
   778 => x"0a",
   779 => x"20",
   780 => x"20",
   781 => x"00",
   782 => x"43",
   783 => x"6d",
   784 => x"64",
   785 => x"5f",
   786 => x"69",
   787 => x"6e",
   788 => x"69",
   789 => x"74",
   790 => x"0a",
   791 => x"00",
   792 => x"43",
   793 => x"4d",
   794 => x"44",
   795 => x"38",
   796 => x"5f",
   797 => x"34",
   798 => x"20",
   799 => x"72",
   800 => x"65",
   801 => x"73",
   802 => x"70",
   803 => x"6f",
   804 => x"6e",
   805 => x"73",
   806 => x"65",
   807 => x"3a",
   808 => x"20",
   809 => x"25",
   810 => x"64",
   811 => x"0a",
   812 => x"00",
   813 => x"43",
   814 => x"4d",
   815 => x"44",
   816 => x"35",
   817 => x"38",
   818 => x"20",
   819 => x"25",
   820 => x"64",
   821 => x"0a",
   822 => x"20",
   823 => x"20",
   824 => x"00",
   825 => x"43",
   826 => x"4d",
   827 => x"44",
   828 => x"35",
   829 => x"38",
   830 => x"5f",
   831 => x"32",
   832 => x"20",
   833 => x"25",
   834 => x"64",
   835 => x"0a",
   836 => x"20",
   837 => x"20",
   838 => x"00",
   839 => x"43",
   840 => x"4d",
   841 => x"44",
   842 => x"35",
   843 => x"38",
   844 => x"20",
   845 => x"25",
   846 => x"64",
   847 => x"0a",
   848 => x"20",
   849 => x"20",
   850 => x"00",
   851 => x"53",
   852 => x"44",
   853 => x"48",
   854 => x"43",
   855 => x"20",
   856 => x"49",
   857 => x"6e",
   858 => x"69",
   859 => x"74",
   860 => x"69",
   861 => x"61",
   862 => x"6c",
   863 => x"69",
   864 => x"7a",
   865 => x"61",
   866 => x"74",
   867 => x"69",
   868 => x"6f",
   869 => x"6e",
   870 => x"20",
   871 => x"65",
   872 => x"72",
   873 => x"72",
   874 => x"6f",
   875 => x"72",
   876 => x"21",
   877 => x"0a",
   878 => x"00",
   879 => x"63",
   880 => x"6d",
   881 => x"64",
   882 => x"5f",
   883 => x"43",
   884 => x"4d",
   885 => x"44",
   886 => x"38",
   887 => x"20",
   888 => x"72",
   889 => x"65",
   890 => x"73",
   891 => x"70",
   892 => x"6f",
   893 => x"6e",
   894 => x"73",
   895 => x"65",
   896 => x"3a",
   897 => x"20",
   898 => x"25",
   899 => x"64",
   900 => x"0a",
   901 => x"00",
   902 => x"52",
   903 => x"65",
   904 => x"61",
   905 => x"64",
   906 => x"20",
   907 => x"63",
   908 => x"6f",
   909 => x"6d",
   910 => x"6d",
   911 => x"61",
   912 => x"6e",
   913 => x"64",
   914 => x"20",
   915 => x"66",
   916 => x"61",
   917 => x"69",
   918 => x"6c",
   919 => x"65",
   920 => x"64",
   921 => x"20",
   922 => x"61",
   923 => x"74",
   924 => x"20",
   925 => x"25",
   926 => x"64",
   927 => x"20",
   928 => x"28",
   929 => x"25",
   930 => x"64",
   931 => x"29",
   932 => x"0a",
   933 => x"00",
   934 => x"1e",
   935 => x"73",
   936 => x"1e",
   937 => x"e1",
   938 => x"48",
   939 => x"c3",
   940 => x"ff",
   941 => x"50",
   942 => x"cc",
   943 => x"ce",
   944 => x"49",
   945 => x"c0",
   946 => x"e4",
   947 => x"da",
   948 => x"87",
   949 => x"d3",
   950 => x"4b",
   951 => x"c0",
   952 => x"1e",
   953 => x"c0",
   954 => x"ff",
   955 => x"f0",
   956 => x"c1",
   957 => x"c1",
   958 => x"49",
   959 => x"f7",
   960 => x"f6",
   961 => x"87",
   962 => x"c4",
   963 => x"86",
   964 => x"70",
   965 => x"98",
   966 => x"05",
   967 => x"c9",
   968 => x"87",
   969 => x"e1",
   970 => x"48",
   971 => x"c3",
   972 => x"ff",
   973 => x"50",
   974 => x"c1",
   975 => x"48",
   976 => x"cb",
   977 => x"87",
   978 => x"fa",
   979 => x"d9",
   980 => x"87",
   981 => x"c1",
   982 => x"8b",
   983 => x"05",
   984 => x"ff",
   985 => x"dc",
   986 => x"87",
   987 => x"c0",
   988 => x"48",
   989 => x"fa",
   990 => x"ca",
   991 => x"87",
   992 => x"1e",
   993 => x"73",
   994 => x"1e",
   995 => x"1e",
   996 => x"fa",
   997 => x"c7",
   998 => x"87",
   999 => x"c6",
  1000 => x"ea",
  1001 => x"1e",
  1002 => x"c0",
  1003 => x"e1",
  1004 => x"f0",
  1005 => x"c1",
  1006 => x"c8",
  1007 => x"49",
  1008 => x"f7",
  1009 => x"c5",
  1010 => x"87",
  1011 => x"70",
  1012 => x"4b",
  1013 => x"73",
  1014 => x"1e",
  1015 => x"cd",
  1016 => x"ef",
  1017 => x"49",
  1018 => x"c0",
  1019 => x"f0",
  1020 => x"e0",
  1021 => x"87",
  1022 => x"c8",
  1023 => x"86",
  1024 => x"c1",
  1025 => x"ab",
  1026 => x"02",
  1027 => x"c8",
  1028 => x"87",
  1029 => x"fe",
  1030 => x"de",
  1031 => x"87",
  1032 => x"c0",
  1033 => x"48",
  1034 => x"c1",
  1035 => x"ff",
  1036 => x"87",
  1037 => x"f5",
  1038 => x"c0",
  1039 => x"87",
  1040 => x"70",
  1041 => x"49",
  1042 => x"cf",
  1043 => x"ff",
  1044 => x"ff",
  1045 => x"99",
  1046 => x"c6",
  1047 => x"ea",
  1048 => x"a9",
  1049 => x"02",
  1050 => x"c8",
  1051 => x"87",
  1052 => x"fe",
  1053 => x"c7",
  1054 => x"87",
  1055 => x"c0",
  1056 => x"48",
  1057 => x"c1",
  1058 => x"e8",
  1059 => x"87",
  1060 => x"e1",
  1061 => x"48",
  1062 => x"c3",
  1063 => x"ff",
  1064 => x"50",
  1065 => x"c0",
  1066 => x"f1",
  1067 => x"4b",
  1068 => x"f9",
  1069 => x"d2",
  1070 => x"87",
  1071 => x"70",
  1072 => x"98",
  1073 => x"02",
  1074 => x"c1",
  1075 => x"c6",
  1076 => x"87",
  1077 => x"c0",
  1078 => x"1e",
  1079 => x"c0",
  1080 => x"ff",
  1081 => x"f0",
  1082 => x"c1",
  1083 => x"fa",
  1084 => x"49",
  1085 => x"f5",
  1086 => x"f8",
  1087 => x"87",
  1088 => x"c4",
  1089 => x"86",
  1090 => x"70",
  1091 => x"98",
  1092 => x"05",
  1093 => x"c0",
  1094 => x"f3",
  1095 => x"87",
  1096 => x"e1",
  1097 => x"48",
  1098 => x"c3",
  1099 => x"ff",
  1100 => x"50",
  1101 => x"e1",
  1102 => x"97",
  1103 => x"bf",
  1104 => x"48",
  1105 => x"c4",
  1106 => x"a6",
  1107 => x"58",
  1108 => x"6e",
  1109 => x"49",
  1110 => x"c3",
  1111 => x"ff",
  1112 => x"99",
  1113 => x"e1",
  1114 => x"48",
  1115 => x"c3",
  1116 => x"ff",
  1117 => x"50",
  1118 => x"e1",
  1119 => x"48",
  1120 => x"c3",
  1121 => x"ff",
  1122 => x"50",
  1123 => x"e1",
  1124 => x"48",
  1125 => x"c3",
  1126 => x"ff",
  1127 => x"50",
  1128 => x"e1",
  1129 => x"48",
  1130 => x"c3",
  1131 => x"ff",
  1132 => x"50",
  1133 => x"c1",
  1134 => x"c0",
  1135 => x"99",
  1136 => x"02",
  1137 => x"c4",
  1138 => x"87",
  1139 => x"c1",
  1140 => x"48",
  1141 => x"d5",
  1142 => x"87",
  1143 => x"c0",
  1144 => x"48",
  1145 => x"d1",
  1146 => x"87",
  1147 => x"c2",
  1148 => x"ab",
  1149 => x"05",
  1150 => x"c4",
  1151 => x"87",
  1152 => x"c0",
  1153 => x"48",
  1154 => x"c8",
  1155 => x"87",
  1156 => x"c1",
  1157 => x"8b",
  1158 => x"05",
  1159 => x"fe",
  1160 => x"e2",
  1161 => x"87",
  1162 => x"c0",
  1163 => x"48",
  1164 => x"26",
  1165 => x"f7",
  1166 => x"da",
  1167 => x"87",
  1168 => x"1e",
  1169 => x"73",
  1170 => x"1e",
  1171 => x"c1",
  1172 => x"c2",
  1173 => x"d8",
  1174 => x"48",
  1175 => x"c1",
  1176 => x"78",
  1177 => x"e9",
  1178 => x"48",
  1179 => x"c3",
  1180 => x"ef",
  1181 => x"50",
  1182 => x"c7",
  1183 => x"4b",
  1184 => x"e5",
  1185 => x"48",
  1186 => x"c3",
  1187 => x"50",
  1188 => x"f7",
  1189 => x"c7",
  1190 => x"87",
  1191 => x"e5",
  1192 => x"48",
  1193 => x"c2",
  1194 => x"50",
  1195 => x"e1",
  1196 => x"48",
  1197 => x"c3",
  1198 => x"ff",
  1199 => x"50",
  1200 => x"c0",
  1201 => x"1e",
  1202 => x"c0",
  1203 => x"e5",
  1204 => x"d0",
  1205 => x"c1",
  1206 => x"c0",
  1207 => x"49",
  1208 => x"f3",
  1209 => x"fd",
  1210 => x"87",
  1211 => x"c4",
  1212 => x"86",
  1213 => x"c1",
  1214 => x"a8",
  1215 => x"05",
  1216 => x"c2",
  1217 => x"87",
  1218 => x"c1",
  1219 => x"4b",
  1220 => x"c2",
  1221 => x"ab",
  1222 => x"05",
  1223 => x"c5",
  1224 => x"87",
  1225 => x"c0",
  1226 => x"48",
  1227 => x"c0",
  1228 => x"f1",
  1229 => x"87",
  1230 => x"c1",
  1231 => x"8b",
  1232 => x"05",
  1233 => x"ff",
  1234 => x"cc",
  1235 => x"87",
  1236 => x"fc",
  1237 => x"c9",
  1238 => x"87",
  1239 => x"c1",
  1240 => x"c2",
  1241 => x"dc",
  1242 => x"58",
  1243 => x"c1",
  1244 => x"c2",
  1245 => x"d8",
  1246 => x"bf",
  1247 => x"05",
  1248 => x"cd",
  1249 => x"87",
  1250 => x"c1",
  1251 => x"1e",
  1252 => x"c0",
  1253 => x"ff",
  1254 => x"f0",
  1255 => x"c1",
  1256 => x"d0",
  1257 => x"49",
  1258 => x"f3",
  1259 => x"cb",
  1260 => x"87",
  1261 => x"c4",
  1262 => x"86",
  1263 => x"e1",
  1264 => x"48",
  1265 => x"c3",
  1266 => x"ff",
  1267 => x"50",
  1268 => x"e5",
  1269 => x"48",
  1270 => x"c3",
  1271 => x"50",
  1272 => x"e1",
  1273 => x"48",
  1274 => x"c3",
  1275 => x"ff",
  1276 => x"50",
  1277 => x"c1",
  1278 => x"48",
  1279 => x"f5",
  1280 => x"e8",
  1281 => x"87",
  1282 => x"0e",
  1283 => x"5e",
  1284 => x"5b",
  1285 => x"5c",
  1286 => x"5d",
  1287 => x"0e",
  1288 => x"1e",
  1289 => x"71",
  1290 => x"4a",
  1291 => x"c0",
  1292 => x"4d",
  1293 => x"e1",
  1294 => x"48",
  1295 => x"c3",
  1296 => x"ff",
  1297 => x"50",
  1298 => x"e5",
  1299 => x"48",
  1300 => x"c2",
  1301 => x"50",
  1302 => x"e9",
  1303 => x"48",
  1304 => x"c7",
  1305 => x"50",
  1306 => x"e1",
  1307 => x"48",
  1308 => x"c3",
  1309 => x"ff",
  1310 => x"50",
  1311 => x"72",
  1312 => x"1e",
  1313 => x"c0",
  1314 => x"ff",
  1315 => x"f0",
  1316 => x"c1",
  1317 => x"d1",
  1318 => x"49",
  1319 => x"f2",
  1320 => x"ce",
  1321 => x"87",
  1322 => x"c4",
  1323 => x"86",
  1324 => x"70",
  1325 => x"98",
  1326 => x"05",
  1327 => x"c1",
  1328 => x"c9",
  1329 => x"87",
  1330 => x"c5",
  1331 => x"ee",
  1332 => x"cd",
  1333 => x"df",
  1334 => x"4b",
  1335 => x"e1",
  1336 => x"48",
  1337 => x"c3",
  1338 => x"ff",
  1339 => x"50",
  1340 => x"e1",
  1341 => x"97",
  1342 => x"bf",
  1343 => x"48",
  1344 => x"c4",
  1345 => x"a6",
  1346 => x"58",
  1347 => x"6e",
  1348 => x"49",
  1349 => x"c3",
  1350 => x"ff",
  1351 => x"99",
  1352 => x"c3",
  1353 => x"fe",
  1354 => x"a9",
  1355 => x"05",
  1356 => x"de",
  1357 => x"87",
  1358 => x"c0",
  1359 => x"4c",
  1360 => x"ef",
  1361 => x"fd",
  1362 => x"87",
  1363 => x"d4",
  1364 => x"66",
  1365 => x"08",
  1366 => x"78",
  1367 => x"08",
  1368 => x"d4",
  1369 => x"66",
  1370 => x"48",
  1371 => x"c4",
  1372 => x"80",
  1373 => x"d8",
  1374 => x"a6",
  1375 => x"58",
  1376 => x"c1",
  1377 => x"84",
  1378 => x"c2",
  1379 => x"c0",
  1380 => x"b7",
  1381 => x"ac",
  1382 => x"04",
  1383 => x"e7",
  1384 => x"87",
  1385 => x"c1",
  1386 => x"4b",
  1387 => x"4d",
  1388 => x"c1",
  1389 => x"8b",
  1390 => x"05",
  1391 => x"ff",
  1392 => x"c5",
  1393 => x"87",
  1394 => x"e1",
  1395 => x"48",
  1396 => x"c3",
  1397 => x"ff",
  1398 => x"50",
  1399 => x"e5",
  1400 => x"48",
  1401 => x"c3",
  1402 => x"50",
  1403 => x"75",
  1404 => x"48",
  1405 => x"26",
  1406 => x"f3",
  1407 => x"e5",
  1408 => x"87",
  1409 => x"1e",
  1410 => x"73",
  1411 => x"1e",
  1412 => x"71",
  1413 => x"4b",
  1414 => x"73",
  1415 => x"49",
  1416 => x"d8",
  1417 => x"29",
  1418 => x"c3",
  1419 => x"ff",
  1420 => x"99",
  1421 => x"73",
  1422 => x"4a",
  1423 => x"c8",
  1424 => x"2a",
  1425 => x"cf",
  1426 => x"fc",
  1427 => x"c0",
  1428 => x"9a",
  1429 => x"72",
  1430 => x"b1",
  1431 => x"73",
  1432 => x"4a",
  1433 => x"c8",
  1434 => x"32",
  1435 => x"c0",
  1436 => x"ff",
  1437 => x"f0",
  1438 => x"c0",
  1439 => x"c0",
  1440 => x"9a",
  1441 => x"72",
  1442 => x"b1",
  1443 => x"73",
  1444 => x"4a",
  1445 => x"d8",
  1446 => x"32",
  1447 => x"ff",
  1448 => x"c0",
  1449 => x"c0",
  1450 => x"c0",
  1451 => x"c0",
  1452 => x"9a",
  1453 => x"72",
  1454 => x"b1",
  1455 => x"71",
  1456 => x"48",
  1457 => x"c4",
  1458 => x"87",
  1459 => x"26",
  1460 => x"4d",
  1461 => x"26",
  1462 => x"4c",
  1463 => x"26",
  1464 => x"4b",
  1465 => x"26",
  1466 => x"4f",
  1467 => x"1e",
  1468 => x"73",
  1469 => x"1e",
  1470 => x"71",
  1471 => x"4b",
  1472 => x"73",
  1473 => x"49",
  1474 => x"c8",
  1475 => x"29",
  1476 => x"c3",
  1477 => x"ff",
  1478 => x"99",
  1479 => x"73",
  1480 => x"4a",
  1481 => x"c8",
  1482 => x"32",
  1483 => x"cf",
  1484 => x"fc",
  1485 => x"c0",
  1486 => x"9a",
  1487 => x"72",
  1488 => x"b1",
  1489 => x"71",
  1490 => x"48",
  1491 => x"e2",
  1492 => x"87",
  1493 => x"0e",
  1494 => x"5e",
  1495 => x"5b",
  1496 => x"5c",
  1497 => x"0e",
  1498 => x"71",
  1499 => x"4b",
  1500 => x"c0",
  1501 => x"4c",
  1502 => x"d0",
  1503 => x"66",
  1504 => x"48",
  1505 => x"c0",
  1506 => x"b7",
  1507 => x"a8",
  1508 => x"06",
  1509 => x"c0",
  1510 => x"e3",
  1511 => x"87",
  1512 => x"13",
  1513 => x"4a",
  1514 => x"cc",
  1515 => x"66",
  1516 => x"97",
  1517 => x"bf",
  1518 => x"49",
  1519 => x"cc",
  1520 => x"66",
  1521 => x"48",
  1522 => x"c1",
  1523 => x"80",
  1524 => x"d0",
  1525 => x"a6",
  1526 => x"58",
  1527 => x"71",
  1528 => x"b7",
  1529 => x"aa",
  1530 => x"02",
  1531 => x"c4",
  1532 => x"87",
  1533 => x"c1",
  1534 => x"48",
  1535 => x"cc",
  1536 => x"87",
  1537 => x"c1",
  1538 => x"84",
  1539 => x"d0",
  1540 => x"66",
  1541 => x"b7",
  1542 => x"ac",
  1543 => x"04",
  1544 => x"ff",
  1545 => x"dd",
  1546 => x"87",
  1547 => x"c0",
  1548 => x"48",
  1549 => x"c2",
  1550 => x"87",
  1551 => x"26",
  1552 => x"4d",
  1553 => x"26",
  1554 => x"4c",
  1555 => x"26",
  1556 => x"4b",
  1557 => x"26",
  1558 => x"4f",
  1559 => x"0e",
  1560 => x"5e",
  1561 => x"5b",
  1562 => x"5c",
  1563 => x"5d",
  1564 => x"0e",
  1565 => x"c1",
  1566 => x"cb",
  1567 => x"da",
  1568 => x"48",
  1569 => x"ff",
  1570 => x"78",
  1571 => x"c1",
  1572 => x"ca",
  1573 => x"ea",
  1574 => x"48",
  1575 => x"c0",
  1576 => x"78",
  1577 => x"c0",
  1578 => x"e6",
  1579 => x"cc",
  1580 => x"49",
  1581 => x"da",
  1582 => x"df",
  1583 => x"87",
  1584 => x"c1",
  1585 => x"c2",
  1586 => x"e2",
  1587 => x"1e",
  1588 => x"c0",
  1589 => x"49",
  1590 => x"fb",
  1591 => x"c9",
  1592 => x"87",
  1593 => x"c4",
  1594 => x"86",
  1595 => x"70",
  1596 => x"98",
  1597 => x"05",
  1598 => x"c5",
  1599 => x"87",
  1600 => x"c0",
  1601 => x"48",
  1602 => x"cb",
  1603 => x"c1",
  1604 => x"87",
  1605 => x"c0",
  1606 => x"4b",
  1607 => x"c1",
  1608 => x"cb",
  1609 => x"d6",
  1610 => x"48",
  1611 => x"c1",
  1612 => x"78",
  1613 => x"c8",
  1614 => x"1e",
  1615 => x"c0",
  1616 => x"e6",
  1617 => x"d9",
  1618 => x"1e",
  1619 => x"c1",
  1620 => x"c3",
  1621 => x"d8",
  1622 => x"49",
  1623 => x"fd",
  1624 => x"fb",
  1625 => x"87",
  1626 => x"c8",
  1627 => x"86",
  1628 => x"70",
  1629 => x"98",
  1630 => x"05",
  1631 => x"c6",
  1632 => x"87",
  1633 => x"c1",
  1634 => x"cb",
  1635 => x"d6",
  1636 => x"48",
  1637 => x"c0",
  1638 => x"78",
  1639 => x"c8",
  1640 => x"1e",
  1641 => x"c0",
  1642 => x"e6",
  1643 => x"e2",
  1644 => x"1e",
  1645 => x"c1",
  1646 => x"c3",
  1647 => x"f4",
  1648 => x"49",
  1649 => x"fd",
  1650 => x"e1",
  1651 => x"87",
  1652 => x"c8",
  1653 => x"86",
  1654 => x"70",
  1655 => x"98",
  1656 => x"05",
  1657 => x"c6",
  1658 => x"87",
  1659 => x"c1",
  1660 => x"cb",
  1661 => x"d6",
  1662 => x"48",
  1663 => x"c0",
  1664 => x"78",
  1665 => x"c8",
  1666 => x"1e",
  1667 => x"c0",
  1668 => x"e6",
  1669 => x"eb",
  1670 => x"1e",
  1671 => x"c1",
  1672 => x"c3",
  1673 => x"f4",
  1674 => x"49",
  1675 => x"fd",
  1676 => x"c7",
  1677 => x"87",
  1678 => x"c8",
  1679 => x"86",
  1680 => x"70",
  1681 => x"98",
  1682 => x"05",
  1683 => x"c5",
  1684 => x"87",
  1685 => x"c0",
  1686 => x"48",
  1687 => x"c9",
  1688 => x"ec",
  1689 => x"87",
  1690 => x"c1",
  1691 => x"cb",
  1692 => x"d6",
  1693 => x"bf",
  1694 => x"1e",
  1695 => x"c0",
  1696 => x"e6",
  1697 => x"f4",
  1698 => x"1e",
  1699 => x"c0",
  1700 => x"e5",
  1701 => x"f7",
  1702 => x"87",
  1703 => x"c8",
  1704 => x"86",
  1705 => x"c1",
  1706 => x"cb",
  1707 => x"d6",
  1708 => x"bf",
  1709 => x"02",
  1710 => x"c1",
  1711 => x"f4",
  1712 => x"87",
  1713 => x"c1",
  1714 => x"c2",
  1715 => x"e2",
  1716 => x"4d",
  1717 => x"48",
  1718 => x"c6",
  1719 => x"fe",
  1720 => x"a0",
  1721 => x"4c",
  1722 => x"c8",
  1723 => x"c0",
  1724 => x"1e",
  1725 => x"70",
  1726 => x"49",
  1727 => x"d8",
  1728 => x"f6",
  1729 => x"87",
  1730 => x"c4",
  1731 => x"86",
  1732 => x"c8",
  1733 => x"a4",
  1734 => x"49",
  1735 => x"69",
  1736 => x"4b",
  1737 => x"c1",
  1738 => x"ca",
  1739 => x"e0",
  1740 => x"9f",
  1741 => x"bf",
  1742 => x"49",
  1743 => x"c5",
  1744 => x"d6",
  1745 => x"ea",
  1746 => x"a9",
  1747 => x"05",
  1748 => x"c0",
  1749 => x"cc",
  1750 => x"87",
  1751 => x"c8",
  1752 => x"a4",
  1753 => x"4a",
  1754 => x"6a",
  1755 => x"49",
  1756 => x"fa",
  1757 => x"e2",
  1758 => x"87",
  1759 => x"70",
  1760 => x"4b",
  1761 => x"db",
  1762 => x"87",
  1763 => x"c7",
  1764 => x"fe",
  1765 => x"a5",
  1766 => x"49",
  1767 => x"9f",
  1768 => x"69",
  1769 => x"49",
  1770 => x"ca",
  1771 => x"e9",
  1772 => x"d5",
  1773 => x"a9",
  1774 => x"02",
  1775 => x"c0",
  1776 => x"cc",
  1777 => x"87",
  1778 => x"c0",
  1779 => x"e4",
  1780 => x"c9",
  1781 => x"49",
  1782 => x"d7",
  1783 => x"d6",
  1784 => x"87",
  1785 => x"c0",
  1786 => x"48",
  1787 => x"c8",
  1788 => x"c8",
  1789 => x"87",
  1790 => x"73",
  1791 => x"1e",
  1792 => x"c0",
  1793 => x"e4",
  1794 => x"e7",
  1795 => x"1e",
  1796 => x"c0",
  1797 => x"e4",
  1798 => x"d6",
  1799 => x"87",
  1800 => x"c1",
  1801 => x"c2",
  1802 => x"e2",
  1803 => x"1e",
  1804 => x"73",
  1805 => x"49",
  1806 => x"f7",
  1807 => x"f1",
  1808 => x"87",
  1809 => x"cc",
  1810 => x"86",
  1811 => x"70",
  1812 => x"98",
  1813 => x"05",
  1814 => x"c0",
  1815 => x"c5",
  1816 => x"87",
  1817 => x"c0",
  1818 => x"48",
  1819 => x"c7",
  1820 => x"e8",
  1821 => x"87",
  1822 => x"c0",
  1823 => x"e4",
  1824 => x"ff",
  1825 => x"49",
  1826 => x"d6",
  1827 => x"ea",
  1828 => x"87",
  1829 => x"c8",
  1830 => x"c0",
  1831 => x"1e",
  1832 => x"c1",
  1833 => x"c2",
  1834 => x"e2",
  1835 => x"49",
  1836 => x"d7",
  1837 => x"c9",
  1838 => x"87",
  1839 => x"c0",
  1840 => x"e7",
  1841 => x"c7",
  1842 => x"1e",
  1843 => x"c0",
  1844 => x"e3",
  1845 => x"e7",
  1846 => x"87",
  1847 => x"c8",
  1848 => x"1e",
  1849 => x"c0",
  1850 => x"e7",
  1851 => x"df",
  1852 => x"1e",
  1853 => x"c1",
  1854 => x"c3",
  1855 => x"f4",
  1856 => x"49",
  1857 => x"fa",
  1858 => x"d1",
  1859 => x"87",
  1860 => x"d0",
  1861 => x"86",
  1862 => x"70",
  1863 => x"98",
  1864 => x"05",
  1865 => x"c0",
  1866 => x"c9",
  1867 => x"87",
  1868 => x"c1",
  1869 => x"ca",
  1870 => x"ea",
  1871 => x"48",
  1872 => x"c1",
  1873 => x"78",
  1874 => x"c0",
  1875 => x"e4",
  1876 => x"87",
  1877 => x"c8",
  1878 => x"1e",
  1879 => x"c0",
  1880 => x"e7",
  1881 => x"e8",
  1882 => x"1e",
  1883 => x"c1",
  1884 => x"c3",
  1885 => x"d8",
  1886 => x"49",
  1887 => x"f9",
  1888 => x"f3",
  1889 => x"87",
  1890 => x"c8",
  1891 => x"86",
  1892 => x"70",
  1893 => x"98",
  1894 => x"02",
  1895 => x"c0",
  1896 => x"cf",
  1897 => x"87",
  1898 => x"c0",
  1899 => x"e5",
  1900 => x"e6",
  1901 => x"1e",
  1902 => x"c0",
  1903 => x"e2",
  1904 => x"ec",
  1905 => x"87",
  1906 => x"c4",
  1907 => x"86",
  1908 => x"c0",
  1909 => x"48",
  1910 => x"c6",
  1911 => x"cd",
  1912 => x"87",
  1913 => x"c1",
  1914 => x"ca",
  1915 => x"e0",
  1916 => x"97",
  1917 => x"bf",
  1918 => x"49",
  1919 => x"c1",
  1920 => x"d5",
  1921 => x"a9",
  1922 => x"05",
  1923 => x"c0",
  1924 => x"cd",
  1925 => x"87",
  1926 => x"c1",
  1927 => x"ca",
  1928 => x"e1",
  1929 => x"97",
  1930 => x"bf",
  1931 => x"49",
  1932 => x"c2",
  1933 => x"ea",
  1934 => x"a9",
  1935 => x"02",
  1936 => x"c0",
  1937 => x"c5",
  1938 => x"87",
  1939 => x"c0",
  1940 => x"48",
  1941 => x"c5",
  1942 => x"ee",
  1943 => x"87",
  1944 => x"c1",
  1945 => x"c2",
  1946 => x"e2",
  1947 => x"97",
  1948 => x"bf",
  1949 => x"49",
  1950 => x"c3",
  1951 => x"e9",
  1952 => x"a9",
  1953 => x"02",
  1954 => x"c0",
  1955 => x"d2",
  1956 => x"87",
  1957 => x"c1",
  1958 => x"c2",
  1959 => x"e2",
  1960 => x"97",
  1961 => x"bf",
  1962 => x"49",
  1963 => x"c3",
  1964 => x"eb",
  1965 => x"a9",
  1966 => x"02",
  1967 => x"c0",
  1968 => x"c5",
  1969 => x"87",
  1970 => x"c0",
  1971 => x"48",
  1972 => x"c5",
  1973 => x"cf",
  1974 => x"87",
  1975 => x"c1",
  1976 => x"c2",
  1977 => x"ed",
  1978 => x"97",
  1979 => x"bf",
  1980 => x"49",
  1981 => x"71",
  1982 => x"99",
  1983 => x"05",
  1984 => x"c0",
  1985 => x"cc",
  1986 => x"87",
  1987 => x"c1",
  1988 => x"c2",
  1989 => x"ee",
  1990 => x"97",
  1991 => x"bf",
  1992 => x"49",
  1993 => x"c2",
  1994 => x"a9",
  1995 => x"02",
  1996 => x"c0",
  1997 => x"c5",
  1998 => x"87",
  1999 => x"c0",
  2000 => x"48",
  2001 => x"c4",
  2002 => x"f2",
  2003 => x"87",
  2004 => x"c1",
  2005 => x"c2",
  2006 => x"ef",
  2007 => x"97",
  2008 => x"bf",
  2009 => x"48",
  2010 => x"c1",
  2011 => x"ca",
  2012 => x"e6",
  2013 => x"58",
  2014 => x"c1",
  2015 => x"ca",
  2016 => x"e2",
  2017 => x"bf",
  2018 => x"48",
  2019 => x"c1",
  2020 => x"88",
  2021 => x"c1",
  2022 => x"ca",
  2023 => x"ea",
  2024 => x"58",
  2025 => x"c1",
  2026 => x"c2",
  2027 => x"f0",
  2028 => x"97",
  2029 => x"bf",
  2030 => x"49",
  2031 => x"73",
  2032 => x"81",
  2033 => x"c1",
  2034 => x"c2",
  2035 => x"f1",
  2036 => x"97",
  2037 => x"bf",
  2038 => x"4a",
  2039 => x"c8",
  2040 => x"32",
  2041 => x"c1",
  2042 => x"ca",
  2043 => x"f6",
  2044 => x"48",
  2045 => x"72",
  2046 => x"a1",
  2047 => x"78",
  2048 => x"c1",
  2049 => x"c2",
  2050 => x"f2",
  2051 => x"97",
  2052 => x"bf",
  2053 => x"48",
  2054 => x"c1",
  2055 => x"cb",
  2056 => x"ce",
  2057 => x"58",
  2058 => x"c1",
  2059 => x"ca",
  2060 => x"ea",
  2061 => x"bf",
  2062 => x"02",
  2063 => x"c2",
  2064 => x"e2",
  2065 => x"87",
  2066 => x"c8",
  2067 => x"1e",
  2068 => x"c0",
  2069 => x"e6",
  2070 => x"c3",
  2071 => x"1e",
  2072 => x"c1",
  2073 => x"c3",
  2074 => x"f4",
  2075 => x"49",
  2076 => x"f6",
  2077 => x"f6",
  2078 => x"87",
  2079 => x"c8",
  2080 => x"86",
  2081 => x"70",
  2082 => x"98",
  2083 => x"02",
  2084 => x"c0",
  2085 => x"c5",
  2086 => x"87",
  2087 => x"c0",
  2088 => x"48",
  2089 => x"c3",
  2090 => x"da",
  2091 => x"87",
  2092 => x"c1",
  2093 => x"ca",
  2094 => x"e2",
  2095 => x"bf",
  2096 => x"48",
  2097 => x"c4",
  2098 => x"30",
  2099 => x"c1",
  2100 => x"cb",
  2101 => x"d2",
  2102 => x"58",
  2103 => x"c1",
  2104 => x"ca",
  2105 => x"e2",
  2106 => x"bf",
  2107 => x"4a",
  2108 => x"c1",
  2109 => x"cb",
  2110 => x"ca",
  2111 => x"5a",
  2112 => x"c1",
  2113 => x"c3",
  2114 => x"c7",
  2115 => x"97",
  2116 => x"bf",
  2117 => x"49",
  2118 => x"c8",
  2119 => x"31",
  2120 => x"c1",
  2121 => x"c3",
  2122 => x"c6",
  2123 => x"97",
  2124 => x"bf",
  2125 => x"4b",
  2126 => x"73",
  2127 => x"a1",
  2128 => x"49",
  2129 => x"c1",
  2130 => x"c3",
  2131 => x"c8",
  2132 => x"97",
  2133 => x"bf",
  2134 => x"4b",
  2135 => x"d0",
  2136 => x"33",
  2137 => x"73",
  2138 => x"a1",
  2139 => x"49",
  2140 => x"c1",
  2141 => x"c3",
  2142 => x"c9",
  2143 => x"97",
  2144 => x"bf",
  2145 => x"4b",
  2146 => x"d8",
  2147 => x"33",
  2148 => x"73",
  2149 => x"a1",
  2150 => x"49",
  2151 => x"c1",
  2152 => x"cb",
  2153 => x"d6",
  2154 => x"59",
  2155 => x"c1",
  2156 => x"cb",
  2157 => x"ca",
  2158 => x"bf",
  2159 => x"91",
  2160 => x"c1",
  2161 => x"ca",
  2162 => x"f6",
  2163 => x"bf",
  2164 => x"81",
  2165 => x"c1",
  2166 => x"ca",
  2167 => x"fe",
  2168 => x"59",
  2169 => x"c1",
  2170 => x"c3",
  2171 => x"cf",
  2172 => x"97",
  2173 => x"bf",
  2174 => x"4b",
  2175 => x"c8",
  2176 => x"33",
  2177 => x"c1",
  2178 => x"c3",
  2179 => x"ce",
  2180 => x"97",
  2181 => x"bf",
  2182 => x"4c",
  2183 => x"74",
  2184 => x"a3",
  2185 => x"4b",
  2186 => x"c1",
  2187 => x"c3",
  2188 => x"d0",
  2189 => x"97",
  2190 => x"bf",
  2191 => x"4c",
  2192 => x"d0",
  2193 => x"34",
  2194 => x"74",
  2195 => x"a3",
  2196 => x"4b",
  2197 => x"c1",
  2198 => x"c3",
  2199 => x"d1",
  2200 => x"97",
  2201 => x"bf",
  2202 => x"4c",
  2203 => x"cf",
  2204 => x"9c",
  2205 => x"d8",
  2206 => x"34",
  2207 => x"74",
  2208 => x"a3",
  2209 => x"4b",
  2210 => x"c1",
  2211 => x"cb",
  2212 => x"c2",
  2213 => x"5b",
  2214 => x"c2",
  2215 => x"8b",
  2216 => x"73",
  2217 => x"92",
  2218 => x"c1",
  2219 => x"cb",
  2220 => x"c2",
  2221 => x"48",
  2222 => x"72",
  2223 => x"a1",
  2224 => x"78",
  2225 => x"c1",
  2226 => x"d0",
  2227 => x"87",
  2228 => x"c1",
  2229 => x"c2",
  2230 => x"f4",
  2231 => x"97",
  2232 => x"bf",
  2233 => x"49",
  2234 => x"c8",
  2235 => x"31",
  2236 => x"c1",
  2237 => x"c2",
  2238 => x"f3",
  2239 => x"97",
  2240 => x"bf",
  2241 => x"4a",
  2242 => x"72",
  2243 => x"a1",
  2244 => x"49",
  2245 => x"c1",
  2246 => x"cb",
  2247 => x"d2",
  2248 => x"59",
  2249 => x"c5",
  2250 => x"31",
  2251 => x"c7",
  2252 => x"ff",
  2253 => x"81",
  2254 => x"c9",
  2255 => x"29",
  2256 => x"c1",
  2257 => x"cb",
  2258 => x"ca",
  2259 => x"59",
  2260 => x"c1",
  2261 => x"c2",
  2262 => x"f9",
  2263 => x"97",
  2264 => x"bf",
  2265 => x"4a",
  2266 => x"c8",
  2267 => x"32",
  2268 => x"c1",
  2269 => x"c2",
  2270 => x"f8",
  2271 => x"97",
  2272 => x"bf",
  2273 => x"4b",
  2274 => x"73",
  2275 => x"a2",
  2276 => x"4a",
  2277 => x"c1",
  2278 => x"cb",
  2279 => x"d6",
  2280 => x"5a",
  2281 => x"c1",
  2282 => x"cb",
  2283 => x"ca",
  2284 => x"bf",
  2285 => x"92",
  2286 => x"c1",
  2287 => x"ca",
  2288 => x"f6",
  2289 => x"bf",
  2290 => x"82",
  2291 => x"c1",
  2292 => x"cb",
  2293 => x"c6",
  2294 => x"5a",
  2295 => x"c1",
  2296 => x"ca",
  2297 => x"fe",
  2298 => x"48",
  2299 => x"c0",
  2300 => x"78",
  2301 => x"c1",
  2302 => x"ca",
  2303 => x"fa",
  2304 => x"48",
  2305 => x"72",
  2306 => x"a1",
  2307 => x"78",
  2308 => x"c1",
  2309 => x"48",
  2310 => x"f4",
  2311 => x"c6",
  2312 => x"87",
  2313 => x"4e",
  2314 => x"6f",
  2315 => x"20",
  2316 => x"70",
  2317 => x"61",
  2318 => x"72",
  2319 => x"74",
  2320 => x"69",
  2321 => x"74",
  2322 => x"69",
  2323 => x"6f",
  2324 => x"6e",
  2325 => x"20",
  2326 => x"73",
  2327 => x"69",
  2328 => x"67",
  2329 => x"6e",
  2330 => x"61",
  2331 => x"74",
  2332 => x"75",
  2333 => x"72",
  2334 => x"65",
  2335 => x"20",
  2336 => x"66",
  2337 => x"6f",
  2338 => x"75",
  2339 => x"6e",
  2340 => x"64",
  2341 => x"0a",
  2342 => x"00",
  2343 => x"52",
  2344 => x"65",
  2345 => x"61",
  2346 => x"64",
  2347 => x"69",
  2348 => x"6e",
  2349 => x"67",
  2350 => x"20",
  2351 => x"62",
  2352 => x"6f",
  2353 => x"6f",
  2354 => x"74",
  2355 => x"20",
  2356 => x"73",
  2357 => x"65",
  2358 => x"63",
  2359 => x"74",
  2360 => x"6f",
  2361 => x"72",
  2362 => x"20",
  2363 => x"25",
  2364 => x"64",
  2365 => x"0a",
  2366 => x"00",
  2367 => x"52",
  2368 => x"65",
  2369 => x"61",
  2370 => x"64",
  2371 => x"20",
  2372 => x"62",
  2373 => x"6f",
  2374 => x"6f",
  2375 => x"74",
  2376 => x"20",
  2377 => x"73",
  2378 => x"65",
  2379 => x"63",
  2380 => x"74",
  2381 => x"6f",
  2382 => x"72",
  2383 => x"20",
  2384 => x"66",
  2385 => x"72",
  2386 => x"6f",
  2387 => x"6d",
  2388 => x"20",
  2389 => x"66",
  2390 => x"69",
  2391 => x"72",
  2392 => x"73",
  2393 => x"74",
  2394 => x"20",
  2395 => x"70",
  2396 => x"61",
  2397 => x"72",
  2398 => x"74",
  2399 => x"69",
  2400 => x"74",
  2401 => x"69",
  2402 => x"6f",
  2403 => x"6e",
  2404 => x"0a",
  2405 => x"00",
  2406 => x"55",
  2407 => x"6e",
  2408 => x"73",
  2409 => x"75",
  2410 => x"70",
  2411 => x"70",
  2412 => x"6f",
  2413 => x"72",
  2414 => x"74",
  2415 => x"65",
  2416 => x"64",
  2417 => x"20",
  2418 => x"70",
  2419 => x"61",
  2420 => x"72",
  2421 => x"74",
  2422 => x"69",
  2423 => x"74",
  2424 => x"69",
  2425 => x"6f",
  2426 => x"6e",
  2427 => x"20",
  2428 => x"74",
  2429 => x"79",
  2430 => x"70",
  2431 => x"65",
  2432 => x"21",
  2433 => x"0d",
  2434 => x"00",
  2435 => x"46",
  2436 => x"41",
  2437 => x"54",
  2438 => x"33",
  2439 => x"32",
  2440 => x"20",
  2441 => x"20",
  2442 => x"20",
  2443 => x"00",
  2444 => x"52",
  2445 => x"65",
  2446 => x"61",
  2447 => x"64",
  2448 => x"69",
  2449 => x"6e",
  2450 => x"67",
  2451 => x"20",
  2452 => x"4d",
  2453 => x"42",
  2454 => x"52",
  2455 => x"0a",
  2456 => x"00",
  2457 => x"46",
  2458 => x"41",
  2459 => x"54",
  2460 => x"31",
  2461 => x"36",
  2462 => x"20",
  2463 => x"20",
  2464 => x"20",
  2465 => x"00",
  2466 => x"46",
  2467 => x"41",
  2468 => x"54",
  2469 => x"33",
  2470 => x"32",
  2471 => x"20",
  2472 => x"20",
  2473 => x"20",
  2474 => x"00",
  2475 => x"46",
  2476 => x"41",
  2477 => x"54",
  2478 => x"31",
  2479 => x"32",
  2480 => x"20",
  2481 => x"20",
  2482 => x"20",
  2483 => x"00",
  2484 => x"50",
  2485 => x"61",
  2486 => x"72",
  2487 => x"74",
  2488 => x"69",
  2489 => x"74",
  2490 => x"69",
  2491 => x"6f",
  2492 => x"6e",
  2493 => x"63",
  2494 => x"6f",
  2495 => x"75",
  2496 => x"6e",
  2497 => x"74",
  2498 => x"20",
  2499 => x"25",
  2500 => x"64",
  2501 => x"0a",
  2502 => x"00",
  2503 => x"48",
  2504 => x"75",
  2505 => x"6e",
  2506 => x"74",
  2507 => x"69",
  2508 => x"6e",
  2509 => x"67",
  2510 => x"20",
  2511 => x"66",
  2512 => x"6f",
  2513 => x"72",
  2514 => x"20",
  2515 => x"66",
  2516 => x"69",
  2517 => x"6c",
  2518 => x"65",
  2519 => x"73",
  2520 => x"79",
  2521 => x"73",
  2522 => x"74",
  2523 => x"65",
  2524 => x"6d",
  2525 => x"0a",
  2526 => x"00",
  2527 => x"46",
  2528 => x"41",
  2529 => x"54",
  2530 => x"33",
  2531 => x"32",
  2532 => x"20",
  2533 => x"20",
  2534 => x"20",
  2535 => x"00",
  2536 => x"46",
  2537 => x"41",
  2538 => x"54",
  2539 => x"31",
  2540 => x"36",
  2541 => x"20",
  2542 => x"20",
  2543 => x"20",
  2544 => x"00",
  2545 => x"52",
  2546 => x"65",
  2547 => x"61",
  2548 => x"64",
  2549 => x"69",
  2550 => x"6e",
  2551 => x"67",
  2552 => x"20",
  2553 => x"64",
  2554 => x"69",
  2555 => x"72",
  2556 => x"65",
  2557 => x"63",
  2558 => x"74",
  2559 => x"6f",
  2560 => x"72",
  2561 => x"79",
  2562 => x"20",
  2563 => x"73",
  2564 => x"65",
  2565 => x"63",
  2566 => x"74",
  2567 => x"6f",
  2568 => x"72",
  2569 => x"20",
  2570 => x"25",
  2571 => x"64",
  2572 => x"0a",
  2573 => x"00",
  2574 => x"66",
  2575 => x"69",
  2576 => x"6c",
  2577 => x"65",
  2578 => x"20",
  2579 => x"22",
  2580 => x"25",
  2581 => x"73",
  2582 => x"22",
  2583 => x"20",
  2584 => x"66",
  2585 => x"6f",
  2586 => x"75",
  2587 => x"6e",
  2588 => x"64",
  2589 => x"0d",
  2590 => x"00",
  2591 => x"47",
  2592 => x"65",
  2593 => x"74",
  2594 => x"46",
  2595 => x"41",
  2596 => x"54",
  2597 => x"4c",
  2598 => x"69",
  2599 => x"6e",
  2600 => x"6b",
  2601 => x"20",
  2602 => x"72",
  2603 => x"65",
  2604 => x"74",
  2605 => x"75",
  2606 => x"72",
  2607 => x"6e",
  2608 => x"65",
  2609 => x"64",
  2610 => x"20",
  2611 => x"25",
  2612 => x"64",
  2613 => x"0a",
  2614 => x"00",
  2615 => x"43",
  2616 => x"61",
  2617 => x"6e",
  2618 => x"27",
  2619 => x"74",
  2620 => x"20",
  2621 => x"6f",
  2622 => x"70",
  2623 => x"65",
  2624 => x"6e",
  2625 => x"20",
  2626 => x"25",
  2627 => x"73",
  2628 => x"0a",
  2629 => x"00",
  2630 => x"0e",
  2631 => x"5e",
  2632 => x"5b",
  2633 => x"5c",
  2634 => x"5d",
  2635 => x"0e",
  2636 => x"71",
  2637 => x"4a",
  2638 => x"c1",
  2639 => x"ca",
  2640 => x"ea",
  2641 => x"bf",
  2642 => x"02",
  2643 => x"cc",
  2644 => x"87",
  2645 => x"72",
  2646 => x"4b",
  2647 => x"c7",
  2648 => x"b7",
  2649 => x"2b",
  2650 => x"72",
  2651 => x"4c",
  2652 => x"c1",
  2653 => x"ff",
  2654 => x"9c",
  2655 => x"ca",
  2656 => x"87",
  2657 => x"72",
  2658 => x"4b",
  2659 => x"c8",
  2660 => x"b7",
  2661 => x"2b",
  2662 => x"72",
  2663 => x"4c",
  2664 => x"c3",
  2665 => x"ff",
  2666 => x"9c",
  2667 => x"c1",
  2668 => x"cb",
  2669 => x"da",
  2670 => x"bf",
  2671 => x"ab",
  2672 => x"02",
  2673 => x"de",
  2674 => x"87",
  2675 => x"c1",
  2676 => x"c2",
  2677 => x"e2",
  2678 => x"1e",
  2679 => x"c1",
  2680 => x"ca",
  2681 => x"f6",
  2682 => x"bf",
  2683 => x"49",
  2684 => x"73",
  2685 => x"81",
  2686 => x"ea",
  2687 => x"c1",
  2688 => x"87",
  2689 => x"c4",
  2690 => x"86",
  2691 => x"70",
  2692 => x"98",
  2693 => x"05",
  2694 => x"c5",
  2695 => x"87",
  2696 => x"c0",
  2697 => x"48",
  2698 => x"c0",
  2699 => x"f6",
  2700 => x"87",
  2701 => x"c1",
  2702 => x"cb",
  2703 => x"de",
  2704 => x"5b",
  2705 => x"c1",
  2706 => x"ca",
  2707 => x"ea",
  2708 => x"bf",
  2709 => x"02",
  2710 => x"d9",
  2711 => x"87",
  2712 => x"74",
  2713 => x"4a",
  2714 => x"c4",
  2715 => x"92",
  2716 => x"c1",
  2717 => x"c2",
  2718 => x"e2",
  2719 => x"82",
  2720 => x"6a",
  2721 => x"49",
  2722 => x"eb",
  2723 => x"dc",
  2724 => x"87",
  2725 => x"70",
  2726 => x"49",
  2727 => x"71",
  2728 => x"4d",
  2729 => x"cf",
  2730 => x"ff",
  2731 => x"ff",
  2732 => x"ff",
  2733 => x"ff",
  2734 => x"9d",
  2735 => x"d0",
  2736 => x"87",
  2737 => x"74",
  2738 => x"4a",
  2739 => x"c2",
  2740 => x"92",
  2741 => x"c1",
  2742 => x"c2",
  2743 => x"e2",
  2744 => x"82",
  2745 => x"9f",
  2746 => x"6a",
  2747 => x"49",
  2748 => x"eb",
  2749 => x"fc",
  2750 => x"87",
  2751 => x"70",
  2752 => x"4d",
  2753 => x"75",
  2754 => x"48",
  2755 => x"ed",
  2756 => x"c9",
  2757 => x"87",
  2758 => x"0e",
  2759 => x"5e",
  2760 => x"5b",
  2761 => x"5c",
  2762 => x"5d",
  2763 => x"0e",
  2764 => x"f4",
  2765 => x"86",
  2766 => x"71",
  2767 => x"4c",
  2768 => x"c0",
  2769 => x"4b",
  2770 => x"c1",
  2771 => x"cb",
  2772 => x"da",
  2773 => x"48",
  2774 => x"ff",
  2775 => x"78",
  2776 => x"c1",
  2777 => x"ca",
  2778 => x"fe",
  2779 => x"bf",
  2780 => x"4d",
  2781 => x"c1",
  2782 => x"cb",
  2783 => x"c2",
  2784 => x"bf",
  2785 => x"7e",
  2786 => x"c1",
  2787 => x"ca",
  2788 => x"ea",
  2789 => x"bf",
  2790 => x"02",
  2791 => x"c9",
  2792 => x"87",
  2793 => x"c1",
  2794 => x"ca",
  2795 => x"e2",
  2796 => x"bf",
  2797 => x"4a",
  2798 => x"c4",
  2799 => x"32",
  2800 => x"c7",
  2801 => x"87",
  2802 => x"c1",
  2803 => x"cb",
  2804 => x"c6",
  2805 => x"bf",
  2806 => x"4a",
  2807 => x"c4",
  2808 => x"32",
  2809 => x"c8",
  2810 => x"a6",
  2811 => x"5a",
  2812 => x"c8",
  2813 => x"a6",
  2814 => x"48",
  2815 => x"c0",
  2816 => x"78",
  2817 => x"c4",
  2818 => x"66",
  2819 => x"48",
  2820 => x"c0",
  2821 => x"a8",
  2822 => x"06",
  2823 => x"c3",
  2824 => x"cf",
  2825 => x"87",
  2826 => x"c8",
  2827 => x"66",
  2828 => x"49",
  2829 => x"cf",
  2830 => x"99",
  2831 => x"05",
  2832 => x"c0",
  2833 => x"e3",
  2834 => x"87",
  2835 => x"6e",
  2836 => x"1e",
  2837 => x"c0",
  2838 => x"e7",
  2839 => x"f1",
  2840 => x"1e",
  2841 => x"d4",
  2842 => x"c2",
  2843 => x"87",
  2844 => x"c1",
  2845 => x"c2",
  2846 => x"e2",
  2847 => x"1e",
  2848 => x"cc",
  2849 => x"66",
  2850 => x"49",
  2851 => x"48",
  2852 => x"c1",
  2853 => x"80",
  2854 => x"d0",
  2855 => x"a6",
  2856 => x"58",
  2857 => x"71",
  2858 => x"49",
  2859 => x"e7",
  2860 => x"d4",
  2861 => x"87",
  2862 => x"cc",
  2863 => x"86",
  2864 => x"c1",
  2865 => x"c2",
  2866 => x"e2",
  2867 => x"4b",
  2868 => x"c3",
  2869 => x"87",
  2870 => x"c0",
  2871 => x"e0",
  2872 => x"83",
  2873 => x"97",
  2874 => x"6b",
  2875 => x"49",
  2876 => x"71",
  2877 => x"99",
  2878 => x"02",
  2879 => x"c2",
  2880 => x"c5",
  2881 => x"87",
  2882 => x"97",
  2883 => x"6b",
  2884 => x"49",
  2885 => x"c3",
  2886 => x"e5",
  2887 => x"a9",
  2888 => x"02",
  2889 => x"c1",
  2890 => x"fb",
  2891 => x"87",
  2892 => x"cb",
  2893 => x"a3",
  2894 => x"49",
  2895 => x"97",
  2896 => x"69",
  2897 => x"49",
  2898 => x"d8",
  2899 => x"99",
  2900 => x"05",
  2901 => x"c1",
  2902 => x"ef",
  2903 => x"87",
  2904 => x"cb",
  2905 => x"1e",
  2906 => x"c0",
  2907 => x"e0",
  2908 => x"66",
  2909 => x"1e",
  2910 => x"73",
  2911 => x"49",
  2912 => x"e9",
  2913 => x"f2",
  2914 => x"87",
  2915 => x"c8",
  2916 => x"86",
  2917 => x"70",
  2918 => x"98",
  2919 => x"05",
  2920 => x"c1",
  2921 => x"dc",
  2922 => x"87",
  2923 => x"dc",
  2924 => x"a3",
  2925 => x"4a",
  2926 => x"6a",
  2927 => x"49",
  2928 => x"e8",
  2929 => x"ce",
  2930 => x"87",
  2931 => x"70",
  2932 => x"4a",
  2933 => x"c4",
  2934 => x"a4",
  2935 => x"49",
  2936 => x"72",
  2937 => x"79",
  2938 => x"da",
  2939 => x"a3",
  2940 => x"4a",
  2941 => x"9f",
  2942 => x"6a",
  2943 => x"49",
  2944 => x"e8",
  2945 => x"f8",
  2946 => x"87",
  2947 => x"c4",
  2948 => x"a6",
  2949 => x"58",
  2950 => x"c1",
  2951 => x"ca",
  2952 => x"ea",
  2953 => x"bf",
  2954 => x"02",
  2955 => x"d8",
  2956 => x"87",
  2957 => x"d4",
  2958 => x"a3",
  2959 => x"4a",
  2960 => x"9f",
  2961 => x"6a",
  2962 => x"49",
  2963 => x"e8",
  2964 => x"e5",
  2965 => x"87",
  2966 => x"70",
  2967 => x"49",
  2968 => x"c0",
  2969 => x"ff",
  2970 => x"ff",
  2971 => x"99",
  2972 => x"71",
  2973 => x"48",
  2974 => x"d0",
  2975 => x"30",
  2976 => x"c8",
  2977 => x"a6",
  2978 => x"58",
  2979 => x"c5",
  2980 => x"87",
  2981 => x"c4",
  2982 => x"a6",
  2983 => x"48",
  2984 => x"c0",
  2985 => x"78",
  2986 => x"c4",
  2987 => x"66",
  2988 => x"4a",
  2989 => x"6e",
  2990 => x"82",
  2991 => x"c8",
  2992 => x"a4",
  2993 => x"49",
  2994 => x"72",
  2995 => x"79",
  2996 => x"c0",
  2997 => x"7c",
  2998 => x"dc",
  2999 => x"66",
  3000 => x"1e",
  3001 => x"c0",
  3002 => x"e8",
  3003 => x"ce",
  3004 => x"1e",
  3005 => x"d1",
  3006 => x"de",
  3007 => x"87",
  3008 => x"c8",
  3009 => x"86",
  3010 => x"c1",
  3011 => x"48",
  3012 => x"c1",
  3013 => x"d0",
  3014 => x"87",
  3015 => x"c8",
  3016 => x"66",
  3017 => x"48",
  3018 => x"c1",
  3019 => x"80",
  3020 => x"cc",
  3021 => x"a6",
  3022 => x"58",
  3023 => x"c8",
  3024 => x"66",
  3025 => x"48",
  3026 => x"c4",
  3027 => x"66",
  3028 => x"a8",
  3029 => x"04",
  3030 => x"fc",
  3031 => x"f1",
  3032 => x"87",
  3033 => x"c1",
  3034 => x"ca",
  3035 => x"ea",
  3036 => x"bf",
  3037 => x"02",
  3038 => x"c0",
  3039 => x"f4",
  3040 => x"87",
  3041 => x"75",
  3042 => x"49",
  3043 => x"f9",
  3044 => x"e0",
  3045 => x"87",
  3046 => x"70",
  3047 => x"4d",
  3048 => x"75",
  3049 => x"1e",
  3050 => x"c0",
  3051 => x"e8",
  3052 => x"df",
  3053 => x"1e",
  3054 => x"d0",
  3055 => x"ed",
  3056 => x"87",
  3057 => x"c8",
  3058 => x"86",
  3059 => x"75",
  3060 => x"49",
  3061 => x"cf",
  3062 => x"ff",
  3063 => x"ff",
  3064 => x"ff",
  3065 => x"f8",
  3066 => x"99",
  3067 => x"a9",
  3068 => x"02",
  3069 => x"d6",
  3070 => x"87",
  3071 => x"75",
  3072 => x"49",
  3073 => x"c2",
  3074 => x"89",
  3075 => x"c1",
  3076 => x"ca",
  3077 => x"e2",
  3078 => x"bf",
  3079 => x"91",
  3080 => x"c1",
  3081 => x"ca",
  3082 => x"fa",
  3083 => x"bf",
  3084 => x"48",
  3085 => x"71",
  3086 => x"80",
  3087 => x"c4",
  3088 => x"a6",
  3089 => x"58",
  3090 => x"fb",
  3091 => x"e7",
  3092 => x"87",
  3093 => x"c0",
  3094 => x"48",
  3095 => x"f4",
  3096 => x"8e",
  3097 => x"e7",
  3098 => x"f3",
  3099 => x"87",
  3100 => x"0e",
  3101 => x"5e",
  3102 => x"5b",
  3103 => x"5c",
  3104 => x"5d",
  3105 => x"0e",
  3106 => x"1e",
  3107 => x"71",
  3108 => x"4b",
  3109 => x"73",
  3110 => x"1e",
  3111 => x"c1",
  3112 => x"cb",
  3113 => x"de",
  3114 => x"49",
  3115 => x"fa",
  3116 => x"d8",
  3117 => x"87",
  3118 => x"c4",
  3119 => x"86",
  3120 => x"70",
  3121 => x"98",
  3122 => x"02",
  3123 => x"c1",
  3124 => x"f7",
  3125 => x"87",
  3126 => x"c1",
  3127 => x"cb",
  3128 => x"e2",
  3129 => x"bf",
  3130 => x"49",
  3131 => x"c7",
  3132 => x"ff",
  3133 => x"81",
  3134 => x"c9",
  3135 => x"29",
  3136 => x"c4",
  3137 => x"a6",
  3138 => x"59",
  3139 => x"c0",
  3140 => x"4d",
  3141 => x"4c",
  3142 => x"6e",
  3143 => x"48",
  3144 => x"c0",
  3145 => x"b7",
  3146 => x"a8",
  3147 => x"06",
  3148 => x"c1",
  3149 => x"ed",
  3150 => x"87",
  3151 => x"c1",
  3152 => x"ca",
  3153 => x"fa",
  3154 => x"bf",
  3155 => x"49",
  3156 => x"c1",
  3157 => x"cb",
  3158 => x"e6",
  3159 => x"bf",
  3160 => x"4a",
  3161 => x"c2",
  3162 => x"8a",
  3163 => x"c1",
  3164 => x"ca",
  3165 => x"e2",
  3166 => x"bf",
  3167 => x"92",
  3168 => x"72",
  3169 => x"a1",
  3170 => x"49",
  3171 => x"c1",
  3172 => x"ca",
  3173 => x"e6",
  3174 => x"bf",
  3175 => x"4a",
  3176 => x"74",
  3177 => x"9a",
  3178 => x"72",
  3179 => x"a1",
  3180 => x"49",
  3181 => x"d4",
  3182 => x"66",
  3183 => x"1e",
  3184 => x"71",
  3185 => x"49",
  3186 => x"e2",
  3187 => x"cd",
  3188 => x"87",
  3189 => x"c4",
  3190 => x"86",
  3191 => x"70",
  3192 => x"98",
  3193 => x"05",
  3194 => x"c5",
  3195 => x"87",
  3196 => x"c0",
  3197 => x"48",
  3198 => x"c1",
  3199 => x"c0",
  3200 => x"87",
  3201 => x"c1",
  3202 => x"84",
  3203 => x"c1",
  3204 => x"ca",
  3205 => x"e6",
  3206 => x"bf",
  3207 => x"49",
  3208 => x"74",
  3209 => x"99",
  3210 => x"05",
  3211 => x"cc",
  3212 => x"87",
  3213 => x"c1",
  3214 => x"cb",
  3215 => x"e6",
  3216 => x"bf",
  3217 => x"49",
  3218 => x"f6",
  3219 => x"f1",
  3220 => x"87",
  3221 => x"c1",
  3222 => x"cb",
  3223 => x"ea",
  3224 => x"58",
  3225 => x"d4",
  3226 => x"66",
  3227 => x"48",
  3228 => x"c8",
  3229 => x"c0",
  3230 => x"80",
  3231 => x"d8",
  3232 => x"a6",
  3233 => x"58",
  3234 => x"c1",
  3235 => x"85",
  3236 => x"6e",
  3237 => x"b7",
  3238 => x"ad",
  3239 => x"04",
  3240 => x"fe",
  3241 => x"e4",
  3242 => x"87",
  3243 => x"cf",
  3244 => x"87",
  3245 => x"73",
  3246 => x"1e",
  3247 => x"c0",
  3248 => x"e8",
  3249 => x"f7",
  3250 => x"1e",
  3251 => x"cd",
  3252 => x"e8",
  3253 => x"87",
  3254 => x"c8",
  3255 => x"86",
  3256 => x"c0",
  3257 => x"48",
  3258 => x"c5",
  3259 => x"87",
  3260 => x"c1",
  3261 => x"cb",
  3262 => x"e2",
  3263 => x"bf",
  3264 => x"48",
  3265 => x"26",
  3266 => x"e5",
  3267 => x"ca",
  3268 => x"87",
  3269 => x"1e",
  3270 => x"f1",
  3271 => x"09",
  3272 => x"97",
  3273 => x"79",
  3274 => x"09",
  3275 => x"71",
  3276 => x"48",
  3277 => x"26",
  3278 => x"4f",
  3279 => x"0e",
  3280 => x"5e",
  3281 => x"5b",
  3282 => x"5c",
  3283 => x"0e",
  3284 => x"71",
  3285 => x"4b",
  3286 => x"c0",
  3287 => x"4c",
  3288 => x"13",
  3289 => x"4a",
  3290 => x"72",
  3291 => x"9a",
  3292 => x"02",
  3293 => x"cd",
  3294 => x"87",
  3295 => x"72",
  3296 => x"49",
  3297 => x"e2",
  3298 => x"87",
  3299 => x"c1",
  3300 => x"84",
  3301 => x"13",
  3302 => x"4a",
  3303 => x"72",
  3304 => x"9a",
  3305 => x"05",
  3306 => x"f3",
  3307 => x"87",
  3308 => x"74",
  3309 => x"48",
  3310 => x"c2",
  3311 => x"87",
  3312 => x"26",
  3313 => x"4d",
  3314 => x"26",
  3315 => x"4c",
  3316 => x"26",
  3317 => x"4b",
  3318 => x"26",
  3319 => x"4f",
  3320 => x"0e",
  3321 => x"5e",
  3322 => x"5b",
  3323 => x"5c",
  3324 => x"5d",
  3325 => x"0e",
  3326 => x"71",
  3327 => x"4b",
  3328 => x"73",
  3329 => x"4c",
  3330 => x"d0",
  3331 => x"66",
  3332 => x"48",
  3333 => x"c2",
  3334 => x"28",
  3335 => x"d4",
  3336 => x"a6",
  3337 => x"58",
  3338 => x"d0",
  3339 => x"66",
  3340 => x"49",
  3341 => x"48",
  3342 => x"c1",
  3343 => x"88",
  3344 => x"d4",
  3345 => x"a6",
  3346 => x"58",
  3347 => x"71",
  3348 => x"99",
  3349 => x"02",
  3350 => x"c1",
  3351 => x"c4",
  3352 => x"87",
  3353 => x"24",
  3354 => x"4d",
  3355 => x"c0",
  3356 => x"4b",
  3357 => x"75",
  3358 => x"4a",
  3359 => x"dc",
  3360 => x"2a",
  3361 => x"c0",
  3362 => x"f0",
  3363 => x"82",
  3364 => x"c0",
  3365 => x"f9",
  3366 => x"aa",
  3367 => x"06",
  3368 => x"c2",
  3369 => x"87",
  3370 => x"c7",
  3371 => x"82",
  3372 => x"72",
  3373 => x"49",
  3374 => x"fe",
  3375 => x"d4",
  3376 => x"87",
  3377 => x"c4",
  3378 => x"35",
  3379 => x"c1",
  3380 => x"83",
  3381 => x"c8",
  3382 => x"b7",
  3383 => x"ab",
  3384 => x"04",
  3385 => x"e2",
  3386 => x"87",
  3387 => x"c0",
  3388 => x"e0",
  3389 => x"49",
  3390 => x"fe",
  3391 => x"c4",
  3392 => x"87",
  3393 => x"d0",
  3394 => x"66",
  3395 => x"49",
  3396 => x"c3",
  3397 => x"99",
  3398 => x"05",
  3399 => x"c5",
  3400 => x"87",
  3401 => x"ca",
  3402 => x"49",
  3403 => x"fd",
  3404 => x"f7",
  3405 => x"87",
  3406 => x"d0",
  3407 => x"66",
  3408 => x"49",
  3409 => x"48",
  3410 => x"c1",
  3411 => x"88",
  3412 => x"d4",
  3413 => x"a6",
  3414 => x"58",
  3415 => x"71",
  3416 => x"99",
  3417 => x"05",
  3418 => x"fe",
  3419 => x"fc",
  3420 => x"87",
  3421 => x"ca",
  3422 => x"49",
  3423 => x"fd",
  3424 => x"e3",
  3425 => x"87",
  3426 => x"26",
  3427 => x"4d",
  3428 => x"26",
  3429 => x"4c",
  3430 => x"26",
  3431 => x"4b",
  3432 => x"26",
  3433 => x"4f",
  3434 => x"0e",
  3435 => x"5e",
  3436 => x"5b",
  3437 => x"5c",
  3438 => x"5d",
  3439 => x"0e",
  3440 => x"fc",
  3441 => x"86",
  3442 => x"71",
  3443 => x"4a",
  3444 => x"c0",
  3445 => x"e0",
  3446 => x"66",
  3447 => x"4c",
  3448 => x"c1",
  3449 => x"cb",
  3450 => x"ea",
  3451 => x"4b",
  3452 => x"c0",
  3453 => x"7e",
  3454 => x"72",
  3455 => x"9a",
  3456 => x"05",
  3457 => x"ce",
  3458 => x"87",
  3459 => x"c1",
  3460 => x"cb",
  3461 => x"eb",
  3462 => x"4b",
  3463 => x"c1",
  3464 => x"cb",
  3465 => x"ea",
  3466 => x"48",
  3467 => x"c0",
  3468 => x"f0",
  3469 => x"50",
  3470 => x"c1",
  3471 => x"d2",
  3472 => x"87",
  3473 => x"72",
  3474 => x"9a",
  3475 => x"02",
  3476 => x"c0",
  3477 => x"e9",
  3478 => x"87",
  3479 => x"d4",
  3480 => x"66",
  3481 => x"4d",
  3482 => x"72",
  3483 => x"1e",
  3484 => x"72",
  3485 => x"49",
  3486 => x"75",
  3487 => x"4a",
  3488 => x"ca",
  3489 => x"cf",
  3490 => x"87",
  3491 => x"26",
  3492 => x"4a",
  3493 => x"c0",
  3494 => x"f8",
  3495 => x"d4",
  3496 => x"81",
  3497 => x"11",
  3498 => x"53",
  3499 => x"71",
  3500 => x"1e",
  3501 => x"72",
  3502 => x"49",
  3503 => x"75",
  3504 => x"4a",
  3505 => x"c9",
  3506 => x"fe",
  3507 => x"87",
  3508 => x"70",
  3509 => x"4a",
  3510 => x"26",
  3511 => x"49",
  3512 => x"c1",
  3513 => x"8c",
  3514 => x"72",
  3515 => x"9a",
  3516 => x"05",
  3517 => x"ff",
  3518 => x"da",
  3519 => x"87",
  3520 => x"c0",
  3521 => x"b7",
  3522 => x"ac",
  3523 => x"06",
  3524 => x"dd",
  3525 => x"87",
  3526 => x"c0",
  3527 => x"e4",
  3528 => x"66",
  3529 => x"02",
  3530 => x"c5",
  3531 => x"87",
  3532 => x"c0",
  3533 => x"f0",
  3534 => x"4a",
  3535 => x"c3",
  3536 => x"87",
  3537 => x"c0",
  3538 => x"e0",
  3539 => x"4a",
  3540 => x"73",
  3541 => x"0a",
  3542 => x"97",
  3543 => x"7a",
  3544 => x"0a",
  3545 => x"c1",
  3546 => x"83",
  3547 => x"8c",
  3548 => x"c0",
  3549 => x"b7",
  3550 => x"ac",
  3551 => x"01",
  3552 => x"ff",
  3553 => x"e3",
  3554 => x"87",
  3555 => x"c1",
  3556 => x"cb",
  3557 => x"ea",
  3558 => x"ab",
  3559 => x"02",
  3560 => x"de",
  3561 => x"87",
  3562 => x"d8",
  3563 => x"66",
  3564 => x"4c",
  3565 => x"dc",
  3566 => x"66",
  3567 => x"1e",
  3568 => x"c1",
  3569 => x"8b",
  3570 => x"97",
  3571 => x"6b",
  3572 => x"49",
  3573 => x"74",
  3574 => x"0f",
  3575 => x"c4",
  3576 => x"86",
  3577 => x"6e",
  3578 => x"48",
  3579 => x"c1",
  3580 => x"80",
  3581 => x"c4",
  3582 => x"a6",
  3583 => x"58",
  3584 => x"c1",
  3585 => x"cb",
  3586 => x"ea",
  3587 => x"ab",
  3588 => x"05",
  3589 => x"ff",
  3590 => x"e5",
  3591 => x"87",
  3592 => x"6e",
  3593 => x"48",
  3594 => x"fc",
  3595 => x"8e",
  3596 => x"26",
  3597 => x"4d",
  3598 => x"26",
  3599 => x"4c",
  3600 => x"26",
  3601 => x"4b",
  3602 => x"26",
  3603 => x"4f",
  3604 => x"30",
  3605 => x"31",
  3606 => x"32",
  3607 => x"33",
  3608 => x"34",
  3609 => x"35",
  3610 => x"36",
  3611 => x"37",
  3612 => x"38",
  3613 => x"39",
  3614 => x"41",
  3615 => x"42",
  3616 => x"43",
  3617 => x"44",
  3618 => x"45",
  3619 => x"46",
  3620 => x"00",
  3621 => x"0e",
  3622 => x"5e",
  3623 => x"5b",
  3624 => x"5c",
  3625 => x"5d",
  3626 => x"0e",
  3627 => x"71",
  3628 => x"4b",
  3629 => x"ff",
  3630 => x"4d",
  3631 => x"13",
  3632 => x"4c",
  3633 => x"74",
  3634 => x"9c",
  3635 => x"02",
  3636 => x"d8",
  3637 => x"87",
  3638 => x"c1",
  3639 => x"85",
  3640 => x"d4",
  3641 => x"66",
  3642 => x"1e",
  3643 => x"74",
  3644 => x"49",
  3645 => x"d4",
  3646 => x"66",
  3647 => x"0f",
  3648 => x"c4",
  3649 => x"86",
  3650 => x"74",
  3651 => x"a8",
  3652 => x"05",
  3653 => x"c7",
  3654 => x"87",
  3655 => x"13",
  3656 => x"4c",
  3657 => x"74",
  3658 => x"9c",
  3659 => x"05",
  3660 => x"e8",
  3661 => x"87",
  3662 => x"75",
  3663 => x"48",
  3664 => x"26",
  3665 => x"4d",
  3666 => x"26",
  3667 => x"4c",
  3668 => x"26",
  3669 => x"4b",
  3670 => x"26",
  3671 => x"4f",
  3672 => x"0e",
  3673 => x"5e",
  3674 => x"5b",
  3675 => x"5c",
  3676 => x"5d",
  3677 => x"0e",
  3678 => x"e8",
  3679 => x"86",
  3680 => x"c4",
  3681 => x"a6",
  3682 => x"59",
  3683 => x"c0",
  3684 => x"e8",
  3685 => x"66",
  3686 => x"4d",
  3687 => x"c0",
  3688 => x"4c",
  3689 => x"c8",
  3690 => x"a6",
  3691 => x"48",
  3692 => x"c0",
  3693 => x"78",
  3694 => x"6e",
  3695 => x"97",
  3696 => x"bf",
  3697 => x"4b",
  3698 => x"6e",
  3699 => x"48",
  3700 => x"c1",
  3701 => x"80",
  3702 => x"c4",
  3703 => x"a6",
  3704 => x"58",
  3705 => x"73",
  3706 => x"9b",
  3707 => x"02",
  3708 => x"c6",
  3709 => x"d3",
  3710 => x"87",
  3711 => x"c8",
  3712 => x"66",
  3713 => x"02",
  3714 => x"c5",
  3715 => x"db",
  3716 => x"87",
  3717 => x"cc",
  3718 => x"a6",
  3719 => x"48",
  3720 => x"c0",
  3721 => x"78",
  3722 => x"fc",
  3723 => x"80",
  3724 => x"c0",
  3725 => x"78",
  3726 => x"73",
  3727 => x"4a",
  3728 => x"c0",
  3729 => x"e0",
  3730 => x"8a",
  3731 => x"02",
  3732 => x"c3",
  3733 => x"c6",
  3734 => x"87",
  3735 => x"c3",
  3736 => x"8a",
  3737 => x"02",
  3738 => x"c3",
  3739 => x"c0",
  3740 => x"87",
  3741 => x"c2",
  3742 => x"8a",
  3743 => x"02",
  3744 => x"c2",
  3745 => x"e8",
  3746 => x"87",
  3747 => x"c2",
  3748 => x"8a",
  3749 => x"02",
  3750 => x"c2",
  3751 => x"f4",
  3752 => x"87",
  3753 => x"c4",
  3754 => x"8a",
  3755 => x"02",
  3756 => x"c2",
  3757 => x"ee",
  3758 => x"87",
  3759 => x"c2",
  3760 => x"8a",
  3761 => x"02",
  3762 => x"c2",
  3763 => x"e8",
  3764 => x"87",
  3765 => x"c3",
  3766 => x"8a",
  3767 => x"02",
  3768 => x"c2",
  3769 => x"ea",
  3770 => x"87",
  3771 => x"d4",
  3772 => x"8a",
  3773 => x"02",
  3774 => x"c0",
  3775 => x"f6",
  3776 => x"87",
  3777 => x"d4",
  3778 => x"8a",
  3779 => x"02",
  3780 => x"c1",
  3781 => x"c0",
  3782 => x"87",
  3783 => x"ca",
  3784 => x"8a",
  3785 => x"02",
  3786 => x"c0",
  3787 => x"f2",
  3788 => x"87",
  3789 => x"c1",
  3790 => x"8a",
  3791 => x"02",
  3792 => x"c1",
  3793 => x"e1",
  3794 => x"87",
  3795 => x"c1",
  3796 => x"8a",
  3797 => x"02",
  3798 => x"df",
  3799 => x"87",
  3800 => x"c8",
  3801 => x"8a",
  3802 => x"02",
  3803 => x"c1",
  3804 => x"ce",
  3805 => x"87",
  3806 => x"c4",
  3807 => x"8a",
  3808 => x"02",
  3809 => x"c0",
  3810 => x"e3",
  3811 => x"87",
  3812 => x"c3",
  3813 => x"8a",
  3814 => x"02",
  3815 => x"c0",
  3816 => x"e5",
  3817 => x"87",
  3818 => x"c2",
  3819 => x"8a",
  3820 => x"02",
  3821 => x"c8",
  3822 => x"87",
  3823 => x"c3",
  3824 => x"8a",
  3825 => x"02",
  3826 => x"d3",
  3827 => x"87",
  3828 => x"c1",
  3829 => x"fa",
  3830 => x"87",
  3831 => x"cc",
  3832 => x"a6",
  3833 => x"48",
  3834 => x"ca",
  3835 => x"78",
  3836 => x"c2",
  3837 => x"d2",
  3838 => x"87",
  3839 => x"cc",
  3840 => x"a6",
  3841 => x"48",
  3842 => x"c2",
  3843 => x"78",
  3844 => x"c2",
  3845 => x"ca",
  3846 => x"87",
  3847 => x"cc",
  3848 => x"a6",
  3849 => x"48",
  3850 => x"d0",
  3851 => x"78",
  3852 => x"c2",
  3853 => x"c2",
  3854 => x"87",
  3855 => x"c0",
  3856 => x"f0",
  3857 => x"66",
  3858 => x"1e",
  3859 => x"c0",
  3860 => x"f0",
  3861 => x"66",
  3862 => x"1e",
  3863 => x"c4",
  3864 => x"85",
  3865 => x"75",
  3866 => x"4a",
  3867 => x"c4",
  3868 => x"8a",
  3869 => x"6a",
  3870 => x"49",
  3871 => x"fc",
  3872 => x"c3",
  3873 => x"87",
  3874 => x"c8",
  3875 => x"86",
  3876 => x"70",
  3877 => x"49",
  3878 => x"71",
  3879 => x"a4",
  3880 => x"4c",
  3881 => x"c1",
  3882 => x"e5",
  3883 => x"87",
  3884 => x"c8",
  3885 => x"a6",
  3886 => x"48",
  3887 => x"c1",
  3888 => x"78",
  3889 => x"c1",
  3890 => x"dd",
  3891 => x"87",
  3892 => x"c0",
  3893 => x"f0",
  3894 => x"66",
  3895 => x"1e",
  3896 => x"c4",
  3897 => x"85",
  3898 => x"75",
  3899 => x"4a",
  3900 => x"c4",
  3901 => x"8a",
  3902 => x"6a",
  3903 => x"49",
  3904 => x"c0",
  3905 => x"f0",
  3906 => x"66",
  3907 => x"0f",
  3908 => x"c4",
  3909 => x"86",
  3910 => x"c1",
  3911 => x"84",
  3912 => x"c1",
  3913 => x"c6",
  3914 => x"87",
  3915 => x"c0",
  3916 => x"f0",
  3917 => x"66",
  3918 => x"1e",
  3919 => x"c0",
  3920 => x"e5",
  3921 => x"49",
  3922 => x"c0",
  3923 => x"f0",
  3924 => x"66",
  3925 => x"0f",
  3926 => x"c4",
  3927 => x"86",
  3928 => x"c1",
  3929 => x"84",
  3930 => x"c0",
  3931 => x"f4",
  3932 => x"87",
  3933 => x"c8",
  3934 => x"a6",
  3935 => x"48",
  3936 => x"c1",
  3937 => x"78",
  3938 => x"c0",
  3939 => x"ec",
  3940 => x"87",
  3941 => x"d0",
  3942 => x"a6",
  3943 => x"48",
  3944 => x"c1",
  3945 => x"78",
  3946 => x"f8",
  3947 => x"80",
  3948 => x"c1",
  3949 => x"78",
  3950 => x"c0",
  3951 => x"e0",
  3952 => x"87",
  3953 => x"c0",
  3954 => x"f0",
  3955 => x"ab",
  3956 => x"06",
  3957 => x"da",
  3958 => x"87",
  3959 => x"c0",
  3960 => x"f9",
  3961 => x"ab",
  3962 => x"03",
  3963 => x"d4",
  3964 => x"87",
  3965 => x"d4",
  3966 => x"66",
  3967 => x"49",
  3968 => x"ca",
  3969 => x"91",
  3970 => x"73",
  3971 => x"4a",
  3972 => x"c0",
  3973 => x"f0",
  3974 => x"8a",
  3975 => x"d4",
  3976 => x"a6",
  3977 => x"48",
  3978 => x"72",
  3979 => x"a1",
  3980 => x"78",
  3981 => x"f4",
  3982 => x"80",
  3983 => x"c1",
  3984 => x"78",
  3985 => x"cc",
  3986 => x"66",
  3987 => x"02",
  3988 => x"c1",
  3989 => x"ea",
  3990 => x"87",
  3991 => x"c4",
  3992 => x"85",
  3993 => x"75",
  3994 => x"49",
  3995 => x"c4",
  3996 => x"89",
  3997 => x"a6",
  3998 => x"48",
  3999 => x"69",
  4000 => x"78",
  4001 => x"c1",
  4002 => x"e4",
  4003 => x"ab",
  4004 => x"05",
  4005 => x"d8",
  4006 => x"87",
  4007 => x"c4",
  4008 => x"66",
  4009 => x"48",
  4010 => x"c0",
  4011 => x"b7",
  4012 => x"a8",
  4013 => x"03",
  4014 => x"cf",
  4015 => x"87",
  4016 => x"c0",
  4017 => x"ed",
  4018 => x"49",
  4019 => x"f4",
  4020 => x"cf",
  4021 => x"87",
  4022 => x"c4",
  4023 => x"66",
  4024 => x"48",
  4025 => x"c0",
  4026 => x"08",
  4027 => x"88",
  4028 => x"c8",
  4029 => x"a6",
  4030 => x"58",
  4031 => x"d0",
  4032 => x"66",
  4033 => x"1e",
  4034 => x"d8",
  4035 => x"66",
  4036 => x"1e",
  4037 => x"c0",
  4038 => x"f8",
  4039 => x"66",
  4040 => x"1e",
  4041 => x"c0",
  4042 => x"f8",
  4043 => x"66",
  4044 => x"1e",
  4045 => x"dc",
  4046 => x"66",
  4047 => x"1e",
  4048 => x"d8",
  4049 => x"66",
  4050 => x"49",
  4051 => x"f6",
  4052 => x"d4",
  4053 => x"87",
  4054 => x"d4",
  4055 => x"86",
  4056 => x"70",
  4057 => x"49",
  4058 => x"71",
  4059 => x"a4",
  4060 => x"4c",
  4061 => x"c0",
  4062 => x"e1",
  4063 => x"87",
  4064 => x"c0",
  4065 => x"e5",
  4066 => x"ab",
  4067 => x"05",
  4068 => x"cf",
  4069 => x"87",
  4070 => x"d0",
  4071 => x"a6",
  4072 => x"48",
  4073 => x"c0",
  4074 => x"78",
  4075 => x"c4",
  4076 => x"80",
  4077 => x"c0",
  4078 => x"78",
  4079 => x"f4",
  4080 => x"80",
  4081 => x"c1",
  4082 => x"78",
  4083 => x"cc",
  4084 => x"87",
  4085 => x"c0",
  4086 => x"f0",
  4087 => x"66",
  4088 => x"1e",
  4089 => x"73",
  4090 => x"49",
  4091 => x"c0",
  4092 => x"f0",
  4093 => x"66",
  4094 => x"0f",
  4095 => x"c4",
  4096 => x"86",
  4097 => x"6e",
  4098 => x"97",
  4099 => x"bf",
  4100 => x"4b",
  4101 => x"6e",
  4102 => x"48",
  4103 => x"c1",
  4104 => x"80",
  4105 => x"c4",
  4106 => x"a6",
  4107 => x"58",
  4108 => x"73",
  4109 => x"9b",
  4110 => x"05",
  4111 => x"f9",
  4112 => x"ed",
  4113 => x"87",
  4114 => x"74",
  4115 => x"48",
  4116 => x"e8",
  4117 => x"8e",
  4118 => x"26",
  4119 => x"4d",
  4120 => x"26",
  4121 => x"4c",
  4122 => x"26",
  4123 => x"4b",
  4124 => x"26",
  4125 => x"4f",
  4126 => x"1e",
  4127 => x"c0",
  4128 => x"1e",
  4129 => x"c0",
  4130 => x"f3",
  4131 => x"c5",
  4132 => x"1e",
  4133 => x"d0",
  4134 => x"a6",
  4135 => x"1e",
  4136 => x"d0",
  4137 => x"66",
  4138 => x"49",
  4139 => x"f8",
  4140 => x"ea",
  4141 => x"87",
  4142 => x"f4",
  4143 => x"8e",
  4144 => x"26",
  4145 => x"4f",
  4146 => x"1e",
  4147 => x"73",
  4148 => x"1e",
  4149 => x"72",
  4150 => x"9a",
  4151 => x"02",
  4152 => x"c0",
  4153 => x"e7",
  4154 => x"87",
  4155 => x"c0",
  4156 => x"48",
  4157 => x"c1",
  4158 => x"4b",
  4159 => x"72",
  4160 => x"a9",
  4161 => x"06",
  4162 => x"d1",
  4163 => x"87",
  4164 => x"72",
  4165 => x"82",
  4166 => x"06",
  4167 => x"c9",
  4168 => x"87",
  4169 => x"73",
  4170 => x"83",
  4171 => x"72",
  4172 => x"a9",
  4173 => x"01",
  4174 => x"f4",
  4175 => x"87",
  4176 => x"c3",
  4177 => x"87",
  4178 => x"c1",
  4179 => x"b2",
  4180 => x"3a",
  4181 => x"72",
  4182 => x"a9",
  4183 => x"03",
  4184 => x"89",
  4185 => x"73",
  4186 => x"80",
  4187 => x"07",
  4188 => x"c1",
  4189 => x"2a",
  4190 => x"2b",
  4191 => x"05",
  4192 => x"f3",
  4193 => x"87",
  4194 => x"26",
  4195 => x"4b",
  4196 => x"26",
  4197 => x"4f",
  4198 => x"1e",
  4199 => x"75",
  4200 => x"1e",
  4201 => x"c4",
  4202 => x"4d",
  4203 => x"71",
  4204 => x"b7",
  4205 => x"a1",
  4206 => x"04",
  4207 => x"ff",
  4208 => x"b9",
  4209 => x"c1",
  4210 => x"81",
  4211 => x"c3",
  4212 => x"bd",
  4213 => x"07",
  4214 => x"72",
  4215 => x"b7",
  4216 => x"a2",
  4217 => x"04",
  4218 => x"ff",
  4219 => x"ba",
  4220 => x"c1",
  4221 => x"82",
  4222 => x"c1",
  4223 => x"bd",
  4224 => x"07",
  4225 => x"fe",
  4226 => x"ee",
  4227 => x"87",
  4228 => x"c1",
  4229 => x"2d",
  4230 => x"04",
  4231 => x"ff",
  4232 => x"b8",
  4233 => x"c1",
  4234 => x"80",
  4235 => x"07",
  4236 => x"2d",
  4237 => x"04",
  4238 => x"ff",
  4239 => x"b9",
  4240 => x"c1",
  4241 => x"81",
  4242 => x"07",
  4243 => x"26",
  4244 => x"4d",
  4245 => x"26",
  4246 => x"4f",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;

