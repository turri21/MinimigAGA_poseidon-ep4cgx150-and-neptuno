library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM-2 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
type ram_type is array (0 to 2 ** (maxAddrBitBRAM-3) - 1) of word_t;

signal ram : ram_type :=
(
     0 => (x"01",x"da",x"87",x"04"),
     1 => (x"dd",x"87",x"0e",x"58"),
     2 => (x"5e",x"59",x"5a",x"0e"),
     3 => (x"27",x"00",x"00",x"00"),
     4 => (x"2c",x"0f",x"26",x"4a"),
     5 => (x"26",x"49",x"26",x"48"),
     6 => (x"ff",x"80",x"26",x"08"),
     7 => (x"4f",x"27",x"00",x"00"),
     8 => (x"00",x"2d",x"4f",x"27"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"4f",x"00",x"fd",x"87"),
    11 => (x"4f",x"c1",x"cb",x"f0"),
    12 => (x"4e",x"c9",x"c0",x"86"),
    13 => (x"c1",x"cb",x"f0",x"49"),
    14 => (x"c1",x"c2",x"cc",x"48"),
    15 => (x"89",x"d0",x"89",x"03"),
    16 => (x"c0",x"40",x"40",x"40"),
    17 => (x"40",x"f6",x"87",x"d0"),
    18 => (x"81",x"05",x"c0",x"50"),
    19 => (x"c1",x"89",x"05",x"f9"),
    20 => (x"87",x"c1",x"c2",x"c9"),
    21 => (x"4d",x"c1",x"c2",x"c9"),
    22 => (x"4c",x"74",x"ad",x"02"),
    23 => (x"c4",x"87",x"24",x"0f"),
    24 => (x"f7",x"87",x"c1",x"c0"),
    25 => (x"87",x"c1",x"c2",x"c9"),
    26 => (x"4d",x"c1",x"c2",x"c9"),
    27 => (x"4c",x"74",x"ad",x"02"),
    28 => (x"c6",x"87",x"c4",x"8c"),
    29 => (x"6c",x"0f",x"f5",x"87"),
    30 => (x"00",x"fd",x"87",x"1e"),
    31 => (x"73",x"1e",x"c2",x"c0"),
    32 => (x"c0",x"4b",x"73",x"0f"),
    33 => (x"c4",x"87",x"26",x"4d"),
    34 => (x"26",x"4c",x"26",x"4b"),
    35 => (x"26",x"4f",x"1e",x"e7"),
    36 => (x"48",x"c0",x"e0",x"50"),
    37 => (x"e7",x"48",x"c0",x"e1"),
    38 => (x"50",x"e7",x"48",x"c0"),
    39 => (x"e0",x"50",x"e7",x"48"),
    40 => (x"c0",x"e1",x"50",x"26"),
    41 => (x"4f",x"1e",x"73",x"1e"),
    42 => (x"e7",x"48",x"c0",x"e0"),
    43 => (x"50",x"e7",x"48",x"c0"),
    44 => (x"e1",x"50",x"c6",x"d0"),
    45 => (x"49",x"c0",x"f1",x"fa"),
    46 => (x"87",x"c0",x"fc",x"c0"),
    47 => (x"4b",x"d1",x"c4",x"87"),
    48 => (x"70",x"98",x"02",x"c1"),
    49 => (x"c8",x"87",x"c0",x"ff"),
    50 => (x"f0",x"4b",x"c5",x"f9"),
    51 => (x"49",x"c0",x"f1",x"e2"),
    52 => (x"87",x"d6",x"f7",x"87"),
    53 => (x"70",x"98",x"02",x"c0"),
    54 => (x"e4",x"87",x"c3",x"f0"),
    55 => (x"4b",x"c2",x"c0",x"c0"),
    56 => (x"1e",x"c4",x"e0",x"49"),
    57 => (x"c0",x"ee",x"d8",x"87"),
    58 => (x"c4",x"86",x"70",x"98"),
    59 => (x"02",x"c6",x"87",x"fe"),
    60 => (x"c9",x"87",x"c0",x"e0"),
    61 => (x"87",x"c4",x"ec",x"49"),
    62 => (x"c0",x"f0",x"f7",x"87"),
    63 => (x"d7",x"87",x"c5",x"c1"),
    64 => (x"49",x"c0",x"f0",x"ee"),
    65 => (x"87",x"c5",x"dd",x"49"),
    66 => (x"c0",x"f0",x"e7",x"87"),
    67 => (x"c7",x"87",x"c6",x"e6"),
    68 => (x"49",x"c0",x"f0",x"de"),
    69 => (x"87",x"73",x"49",x"fd"),
    70 => (x"f4",x"87",x"fe",x"d5"),
    71 => (x"87",x"fd",x"ea",x"87"),
    72 => (x"38",x"33",x"32",x"4f"),
    73 => (x"53",x"44",x"41",x"42"),
    74 => (x"42",x"49",x"4e",x"00"),
    75 => (x"43",x"61",x"6e",x"27"),
    76 => (x"74",x"20",x"6c",x"6f"),
    77 => (x"61",x"64",x"20",x"66"),
    78 => (x"69",x"72",x"6d",x"77"),
    79 => (x"61",x"72",x"65",x"0a"),
    80 => (x"00",x"55",x"6e",x"61"),
    81 => (x"62",x"6c",x"65",x"20"),
    82 => (x"74",x"6f",x"20",x"6c"),
    83 => (x"6f",x"63",x"61",x"74"),
    84 => (x"65",x"20",x"70",x"61"),
    85 => (x"72",x"74",x"69",x"74"),
    86 => (x"69",x"6f",x"6e",x"0a"),
    87 => (x"00",x"55",x"6e",x"61"),
    88 => (x"62",x"6c",x"65",x"20"),
    89 => (x"74",x"6f",x"20",x"6c"),
    90 => (x"6f",x"63",x"61",x"74"),
    91 => (x"65",x"20",x"70",x"61"),
    92 => (x"72",x"74",x"69",x"74"),
    93 => (x"69",x"6f",x"6e",x"0a"),
    94 => (x"00",x"48",x"75",x"6e"),
    95 => (x"74",x"69",x"6e",x"67"),
    96 => (x"20",x"66",x"6f",x"72"),
    97 => (x"20",x"70",x"61",x"72"),
    98 => (x"74",x"69",x"74",x"69"),
    99 => (x"6f",x"6e",x"0a",x"00"),
   100 => (x"49",x"6e",x"69",x"74"),
   101 => (x"69",x"61",x"6c",x"69"),
   102 => (x"7a",x"69",x"6e",x"67"),
   103 => (x"20",x"53",x"44",x"20"),
   104 => (x"63",x"61",x"72",x"64"),
   105 => (x"0a",x"00",x"46",x"61"),
   106 => (x"69",x"6c",x"65",x"64"),
   107 => (x"20",x"74",x"6f",x"20"),
   108 => (x"69",x"6e",x"69",x"74"),
   109 => (x"69",x"61",x"6c",x"69"),
   110 => (x"7a",x"65",x"20",x"53"),
   111 => (x"44",x"20",x"63",x"61"),
   112 => (x"72",x"64",x"0a",x"00"),
   113 => (x"1e",x"e4",x"86",x"e3"),
   114 => (x"48",x"c3",x"ff",x"50"),
   115 => (x"e3",x"97",x"bf",x"48"),
   116 => (x"c4",x"a6",x"58",x"6e"),
   117 => (x"49",x"c3",x"ff",x"99"),
   118 => (x"e3",x"48",x"c3",x"ff"),
   119 => (x"50",x"c8",x"31",x"e3"),
   120 => (x"97",x"bf",x"48",x"c8"),
   121 => (x"a6",x"58",x"c4",x"66"),
   122 => (x"48",x"c3",x"ff",x"98"),
   123 => (x"cc",x"a6",x"58",x"c8"),
   124 => (x"66",x"b1",x"e3",x"48"),
   125 => (x"c3",x"ff",x"50",x"c8"),
   126 => (x"31",x"e3",x"97",x"bf"),
   127 => (x"48",x"d0",x"a6",x"58"),
   128 => (x"cc",x"66",x"48",x"c3"),
   129 => (x"ff",x"98",x"d4",x"a6"),
   130 => (x"58",x"d0",x"66",x"b1"),
   131 => (x"e3",x"48",x"c3",x"ff"),
   132 => (x"50",x"c8",x"31",x"e3"),
   133 => (x"97",x"bf",x"48",x"d8"),
   134 => (x"a6",x"58",x"d4",x"66"),
   135 => (x"48",x"c3",x"ff",x"98"),
   136 => (x"dc",x"a6",x"58",x"d8"),
   137 => (x"66",x"b1",x"71",x"48"),
   138 => (x"e4",x"8e",x"26",x"4f"),
   139 => (x"0e",x"5e",x"5b",x"5c"),
   140 => (x"0e",x"1e",x"71",x"4a"),
   141 => (x"72",x"49",x"c3",x"ff"),
   142 => (x"99",x"e3",x"09",x"97"),
   143 => (x"79",x"09",x"c1",x"c2"),
   144 => (x"cc",x"bf",x"05",x"c8"),
   145 => (x"87",x"d0",x"66",x"48"),
   146 => (x"c9",x"30",x"d4",x"a6"),
   147 => (x"58",x"d0",x"66",x"49"),
   148 => (x"d8",x"29",x"c3",x"ff"),
   149 => (x"99",x"e3",x"09",x"97"),
   150 => (x"79",x"09",x"d0",x"66"),
   151 => (x"49",x"d0",x"29",x"c3"),
   152 => (x"ff",x"99",x"e3",x"09"),
   153 => (x"97",x"79",x"09",x"d0"),
   154 => (x"66",x"49",x"c8",x"29"),
   155 => (x"c3",x"ff",x"99",x"e3"),
   156 => (x"09",x"97",x"79",x"09"),
   157 => (x"d0",x"66",x"49",x"c3"),
   158 => (x"ff",x"99",x"e3",x"09"),
   159 => (x"97",x"79",x"09",x"72"),
   160 => (x"49",x"d0",x"29",x"c3"),
   161 => (x"ff",x"99",x"e3",x"09"),
   162 => (x"97",x"79",x"09",x"97"),
   163 => (x"bf",x"48",x"c4",x"a6"),
   164 => (x"58",x"6e",x"4b",x"c3"),
   165 => (x"ff",x"9b",x"c9",x"f0"),
   166 => (x"ff",x"4c",x"c3",x"ff"),
   167 => (x"ab",x"05",x"dc",x"87"),
   168 => (x"e3",x"48",x"c3",x"ff"),
   169 => (x"50",x"e3",x"97",x"bf"),
   170 => (x"48",x"c4",x"a6",x"58"),
   171 => (x"6e",x"4b",x"c3",x"ff"),
   172 => (x"9b",x"c1",x"8c",x"02"),
   173 => (x"c6",x"87",x"c3",x"ff"),
   174 => (x"ab",x"02",x"e4",x"87"),
   175 => (x"73",x"4a",x"c4",x"b7"),
   176 => (x"2a",x"c0",x"f0",x"a2"),
   177 => (x"49",x"c0",x"e9",x"e0"),
   178 => (x"87",x"73",x"4a",x"cf"),
   179 => (x"9a",x"c0",x"f0",x"a2"),
   180 => (x"49",x"c0",x"e9",x"d4"),
   181 => (x"87",x"73",x"48",x"26"),
   182 => (x"c2",x"87",x"26",x"4d"),
   183 => (x"26",x"4c",x"26",x"4b"),
   184 => (x"26",x"4f",x"1e",x"c0"),
   185 => (x"49",x"e3",x"48",x"c3"),
   186 => (x"ff",x"50",x"c1",x"81"),
   187 => (x"c3",x"c8",x"b7",x"a9"),
   188 => (x"04",x"f2",x"87",x"26"),
   189 => (x"4f",x"1e",x"73",x"1e"),
   190 => (x"e8",x"87",x"c4",x"f8"),
   191 => (x"df",x"4b",x"c0",x"1e"),
   192 => (x"c0",x"ff",x"f0",x"c1"),
   193 => (x"f7",x"49",x"fc",x"e3"),
   194 => (x"87",x"c4",x"86",x"c1"),
   195 => (x"a8",x"05",x"c0",x"e8"),
   196 => (x"87",x"e3",x"48",x"c3"),
   197 => (x"ff",x"50",x"c1",x"c0"),
   198 => (x"c0",x"c0",x"c0",x"c0"),
   199 => (x"1e",x"c0",x"e1",x"f0"),
   200 => (x"c1",x"e9",x"49",x"fc"),
   201 => (x"c6",x"87",x"c4",x"86"),
   202 => (x"70",x"98",x"05",x"c9"),
   203 => (x"87",x"e3",x"48",x"c3"),
   204 => (x"ff",x"50",x"c1",x"48"),
   205 => (x"cb",x"87",x"fe",x"e9"),
   206 => (x"87",x"c1",x"8b",x"05"),
   207 => (x"fe",x"ff",x"87",x"c0"),
   208 => (x"48",x"fe",x"da",x"87"),
   209 => (x"43",x"4d",x"44",x"34"),
   210 => (x"31",x"20",x"25",x"64"),
   211 => (x"0a",x"00",x"43",x"4d"),
   212 => (x"44",x"35",x"35",x"20"),
   213 => (x"25",x"64",x"0a",x"00"),
   214 => (x"43",x"4d",x"44",x"34"),
   215 => (x"31",x"20",x"25",x"64"),
   216 => (x"0a",x"00",x"43",x"4d"),
   217 => (x"44",x"35",x"35",x"20"),
   218 => (x"25",x"64",x"0a",x"00"),
   219 => (x"69",x"6e",x"69",x"74"),
   220 => (x"20",x"25",x"64",x"0a"),
   221 => (x"20",x"20",x"00",x"69"),
   222 => (x"6e",x"69",x"74",x"20"),
   223 => (x"25",x"64",x"0a",x"20"),
   224 => (x"20",x"00",x"43",x"6d"),
   225 => (x"64",x"5f",x"69",x"6e"),
   226 => (x"69",x"74",x"0a",x"00"),
   227 => (x"43",x"4d",x"44",x"38"),
   228 => (x"5f",x"34",x"20",x"72"),
   229 => (x"65",x"73",x"70",x"6f"),
   230 => (x"6e",x"73",x"65",x"3a"),
   231 => (x"20",x"25",x"64",x"0a"),
   232 => (x"00",x"43",x"4d",x"44"),
   233 => (x"35",x"38",x"20",x"25"),
   234 => (x"64",x"0a",x"20",x"20"),
   235 => (x"00",x"43",x"4d",x"44"),
   236 => (x"35",x"38",x"5f",x"32"),
   237 => (x"20",x"25",x"64",x"0a"),
   238 => (x"20",x"20",x"00",x"43"),
   239 => (x"4d",x"44",x"35",x"38"),
   240 => (x"20",x"25",x"64",x"0a"),
   241 => (x"20",x"20",x"00",x"53"),
   242 => (x"44",x"48",x"43",x"20"),
   243 => (x"49",x"6e",x"69",x"74"),
   244 => (x"69",x"61",x"6c",x"69"),
   245 => (x"7a",x"61",x"74",x"69"),
   246 => (x"6f",x"6e",x"20",x"65"),
   247 => (x"72",x"72",x"6f",x"72"),
   248 => (x"21",x"0a",x"00",x"63"),
   249 => (x"6d",x"64",x"5f",x"43"),
   250 => (x"4d",x"44",x"38",x"20"),
   251 => (x"72",x"65",x"73",x"70"),
   252 => (x"6f",x"6e",x"73",x"65"),
   253 => (x"3a",x"20",x"25",x"64"),
   254 => (x"0a",x"00",x"52",x"65"),
   255 => (x"61",x"64",x"20",x"63"),
   256 => (x"6f",x"6d",x"6d",x"61"),
   257 => (x"6e",x"64",x"20",x"66"),
   258 => (x"61",x"69",x"6c",x"65"),
   259 => (x"64",x"20",x"61",x"74"),
   260 => (x"20",x"25",x"64",x"20"),
   261 => (x"28",x"25",x"64",x"29"),
   262 => (x"0a",x"00",x"1e",x"73"),
   263 => (x"1e",x"e3",x"48",x"c3"),
   264 => (x"ff",x"50",x"ce",x"c2"),
   265 => (x"49",x"c0",x"e4",x"ca"),
   266 => (x"87",x"d3",x"4b",x"c0"),
   267 => (x"1e",x"c0",x"ff",x"f0"),
   268 => (x"c1",x"c1",x"49",x"f7"),
   269 => (x"f6",x"87",x"c4",x"86"),
   270 => (x"70",x"98",x"05",x"c9"),
   271 => (x"87",x"e3",x"48",x"c3"),
   272 => (x"ff",x"50",x"c1",x"48"),
   273 => (x"cb",x"87",x"fa",x"d9"),
   274 => (x"87",x"c1",x"8b",x"05"),
   275 => (x"ff",x"dc",x"87",x"c0"),
   276 => (x"48",x"fa",x"ca",x"87"),
   277 => (x"1e",x"73",x"1e",x"1e"),
   278 => (x"fa",x"c7",x"87",x"c6"),
   279 => (x"ea",x"1e",x"c0",x"e1"),
   280 => (x"f0",x"c1",x"c8",x"49"),
   281 => (x"f7",x"c5",x"87",x"70"),
   282 => (x"4b",x"73",x"1e",x"cf"),
   283 => (x"e3",x"49",x"c0",x"ee"),
   284 => (x"de",x"87",x"c8",x"86"),
   285 => (x"c1",x"ab",x"02",x"c8"),
   286 => (x"87",x"fe",x"de",x"87"),
   287 => (x"c0",x"48",x"c1",x"ff"),
   288 => (x"87",x"f5",x"c0",x"87"),
   289 => (x"70",x"49",x"cf",x"ff"),
   290 => (x"ff",x"99",x"c6",x"ea"),
   291 => (x"a9",x"02",x"c8",x"87"),
   292 => (x"fe",x"c7",x"87",x"c0"),
   293 => (x"48",x"c1",x"e8",x"87"),
   294 => (x"e3",x"48",x"c3",x"ff"),
   295 => (x"50",x"c0",x"f1",x"4b"),
   296 => (x"f9",x"d2",x"87",x"70"),
   297 => (x"98",x"02",x"c1",x"c6"),
   298 => (x"87",x"c0",x"1e",x"c0"),
   299 => (x"ff",x"f0",x"c1",x"fa"),
   300 => (x"49",x"f5",x"f8",x"87"),
   301 => (x"c4",x"86",x"70",x"98"),
   302 => (x"05",x"c0",x"f3",x"87"),
   303 => (x"e3",x"48",x"c3",x"ff"),
   304 => (x"50",x"e3",x"97",x"bf"),
   305 => (x"48",x"c4",x"a6",x"58"),
   306 => (x"6e",x"49",x"c3",x"ff"),
   307 => (x"99",x"e3",x"48",x"c3"),
   308 => (x"ff",x"50",x"e3",x"48"),
   309 => (x"c3",x"ff",x"50",x"e3"),
   310 => (x"48",x"c3",x"ff",x"50"),
   311 => (x"e3",x"48",x"c3",x"ff"),
   312 => (x"50",x"c1",x"c0",x"99"),
   313 => (x"02",x"c4",x"87",x"c1"),
   314 => (x"48",x"d5",x"87",x"c0"),
   315 => (x"48",x"d1",x"87",x"c2"),
   316 => (x"ab",x"05",x"c4",x"87"),
   317 => (x"c0",x"48",x"c8",x"87"),
   318 => (x"c1",x"8b",x"05",x"fe"),
   319 => (x"e2",x"87",x"c0",x"48"),
   320 => (x"26",x"f7",x"da",x"87"),
   321 => (x"1e",x"73",x"1e",x"c1"),
   322 => (x"c2",x"cc",x"48",x"c1"),
   323 => (x"78",x"eb",x"48",x"c3"),
   324 => (x"ef",x"50",x"c7",x"4b"),
   325 => (x"e7",x"48",x"c3",x"50"),
   326 => (x"f7",x"c7",x"87",x"e7"),
   327 => (x"48",x"c2",x"50",x"e3"),
   328 => (x"48",x"c3",x"ff",x"50"),
   329 => (x"c0",x"1e",x"c0",x"e5"),
   330 => (x"d0",x"c1",x"c0",x"49"),
   331 => (x"f3",x"fd",x"87",x"c4"),
   332 => (x"86",x"c1",x"a8",x"05"),
   333 => (x"c2",x"87",x"c1",x"4b"),
   334 => (x"c2",x"ab",x"05",x"c5"),
   335 => (x"87",x"c0",x"48",x"c0"),
   336 => (x"f1",x"87",x"c1",x"8b"),
   337 => (x"05",x"ff",x"cc",x"87"),
   338 => (x"fc",x"c9",x"87",x"c1"),
   339 => (x"c2",x"d0",x"58",x"c1"),
   340 => (x"c2",x"cc",x"bf",x"05"),
   341 => (x"cd",x"87",x"c1",x"1e"),
   342 => (x"c0",x"ff",x"f0",x"c1"),
   343 => (x"d0",x"49",x"f3",x"cb"),
   344 => (x"87",x"c4",x"86",x"e3"),
   345 => (x"48",x"c3",x"ff",x"50"),
   346 => (x"e7",x"48",x"c3",x"50"),
   347 => (x"e3",x"48",x"c3",x"ff"),
   348 => (x"50",x"c1",x"48",x"f5"),
   349 => (x"e8",x"87",x"0e",x"5e"),
   350 => (x"5b",x"5c",x"5d",x"0e"),
   351 => (x"1e",x"71",x"4a",x"c0"),
   352 => (x"4d",x"e3",x"48",x"c3"),
   353 => (x"ff",x"50",x"e7",x"48"),
   354 => (x"c2",x"50",x"eb",x"48"),
   355 => (x"c7",x"50",x"e3",x"48"),
   356 => (x"c3",x"ff",x"50",x"72"),
   357 => (x"1e",x"c0",x"ff",x"f0"),
   358 => (x"c1",x"d1",x"49",x"f2"),
   359 => (x"ce",x"87",x"c4",x"86"),
   360 => (x"70",x"98",x"05",x"c1"),
   361 => (x"c9",x"87",x"c5",x"ee"),
   362 => (x"cd",x"df",x"4b",x"e3"),
   363 => (x"48",x"c3",x"ff",x"50"),
   364 => (x"e3",x"97",x"bf",x"48"),
   365 => (x"c4",x"a6",x"58",x"6e"),
   366 => (x"49",x"c3",x"ff",x"99"),
   367 => (x"c3",x"fe",x"a9",x"05"),
   368 => (x"de",x"87",x"c0",x"4c"),
   369 => (x"ef",x"fd",x"87",x"d4"),
   370 => (x"66",x"08",x"78",x"08"),
   371 => (x"d4",x"66",x"48",x"c4"),
   372 => (x"80",x"d8",x"a6",x"58"),
   373 => (x"c1",x"84",x"c2",x"c0"),
   374 => (x"b7",x"ac",x"04",x"e7"),
   375 => (x"87",x"c1",x"4b",x"4d"),
   376 => (x"c1",x"8b",x"05",x"ff"),
   377 => (x"c5",x"87",x"e3",x"48"),
   378 => (x"c3",x"ff",x"50",x"e7"),
   379 => (x"48",x"c3",x"50",x"75"),
   380 => (x"48",x"26",x"f3",x"e5"),
   381 => (x"87",x"1e",x"73",x"1e"),
   382 => (x"71",x"4b",x"73",x"49"),
   383 => (x"d8",x"29",x"c3",x"ff"),
   384 => (x"99",x"73",x"4a",x"c8"),
   385 => (x"2a",x"cf",x"fc",x"c0"),
   386 => (x"9a",x"72",x"b1",x"73"),
   387 => (x"4a",x"c8",x"32",x"c0"),
   388 => (x"ff",x"f0",x"c0",x"c0"),
   389 => (x"9a",x"72",x"b1",x"73"),
   390 => (x"4a",x"d8",x"32",x"ff"),
   391 => (x"c0",x"c0",x"c0",x"c0"),
   392 => (x"9a",x"72",x"b1",x"71"),
   393 => (x"48",x"c4",x"87",x"26"),
   394 => (x"4d",x"26",x"4c",x"26"),
   395 => (x"4b",x"26",x"4f",x"1e"),
   396 => (x"73",x"1e",x"71",x"4b"),
   397 => (x"73",x"49",x"c8",x"29"),
   398 => (x"c3",x"ff",x"99",x"73"),
   399 => (x"4a",x"c8",x"32",x"cf"),
   400 => (x"fc",x"c0",x"9a",x"72"),
   401 => (x"b1",x"71",x"48",x"e2"),
   402 => (x"87",x"0e",x"5e",x"5b"),
   403 => (x"5c",x"0e",x"71",x"4b"),
   404 => (x"c0",x"4c",x"d0",x"66"),
   405 => (x"48",x"c0",x"b7",x"a8"),
   406 => (x"06",x"c0",x"e3",x"87"),
   407 => (x"13",x"4a",x"cc",x"66"),
   408 => (x"97",x"bf",x"49",x"cc"),
   409 => (x"66",x"48",x"c1",x"80"),
   410 => (x"d0",x"a6",x"58",x"71"),
   411 => (x"b7",x"aa",x"02",x"c4"),
   412 => (x"87",x"c1",x"48",x"cc"),
   413 => (x"87",x"c1",x"84",x"d0"),
   414 => (x"66",x"b7",x"ac",x"04"),
   415 => (x"ff",x"dd",x"87",x"c0"),
   416 => (x"48",x"c2",x"87",x"26"),
   417 => (x"4d",x"26",x"4c",x"26"),
   418 => (x"4b",x"26",x"4f",x"0e"),
   419 => (x"5e",x"5b",x"5c",x"0e"),
   420 => (x"1e",x"c1",x"cb",x"ce"),
   421 => (x"48",x"ff",x"78",x"c1"),
   422 => (x"ca",x"de",x"48",x"c0"),
   423 => (x"78",x"c0",x"e7",x"f0"),
   424 => (x"49",x"da",x"cf",x"87"),
   425 => (x"c1",x"c2",x"d6",x"1e"),
   426 => (x"c0",x"49",x"fb",x"c9"),
   427 => (x"87",x"c4",x"86",x"70"),
   428 => (x"98",x"05",x"c5",x"87"),
   429 => (x"c0",x"48",x"ca",x"f0"),
   430 => (x"87",x"c0",x"4b",x"c1"),
   431 => (x"cb",x"ca",x"48",x"c1"),
   432 => (x"78",x"c8",x"1e",x"c0"),
   433 => (x"e7",x"fd",x"1e",x"c1"),
   434 => (x"c3",x"cc",x"49",x"fd"),
   435 => (x"fb",x"87",x"c8",x"86"),
   436 => (x"70",x"98",x"05",x"c6"),
   437 => (x"87",x"c1",x"cb",x"ca"),
   438 => (x"48",x"c0",x"78",x"c8"),
   439 => (x"1e",x"c0",x"e8",x"c6"),
   440 => (x"1e",x"c1",x"c3",x"e8"),
   441 => (x"49",x"fd",x"e1",x"87"),
   442 => (x"c8",x"86",x"70",x"98"),
   443 => (x"05",x"c6",x"87",x"c1"),
   444 => (x"cb",x"ca",x"48",x"c0"),
   445 => (x"78",x"c8",x"1e",x"c0"),
   446 => (x"e8",x"cf",x"1e",x"c1"),
   447 => (x"c3",x"e8",x"49",x"fd"),
   448 => (x"c7",x"87",x"c8",x"86"),
   449 => (x"70",x"98",x"05",x"c5"),
   450 => (x"87",x"c0",x"48",x"c9"),
   451 => (x"db",x"87",x"c1",x"cb"),
   452 => (x"ca",x"bf",x"1e",x"c0"),
   453 => (x"e8",x"d8",x"1e",x"c0"),
   454 => (x"e3",x"f5",x"87",x"c8"),
   455 => (x"86",x"c1",x"cb",x"ca"),
   456 => (x"bf",x"02",x"c1",x"ed"),
   457 => (x"87",x"c1",x"c2",x"d6"),
   458 => (x"4a",x"48",x"c6",x"fe"),
   459 => (x"a0",x"4c",x"c1",x"c9"),
   460 => (x"dc",x"bf",x"4b",x"c1"),
   461 => (x"ca",x"d4",x"9f",x"bf"),
   462 => (x"49",x"c4",x"a6",x"5a"),
   463 => (x"c5",x"d6",x"ea",x"a9"),
   464 => (x"05",x"c0",x"cc",x"87"),
   465 => (x"c8",x"a4",x"4a",x"6a"),
   466 => (x"49",x"fa",x"e9",x"87"),
   467 => (x"70",x"4b",x"db",x"87"),
   468 => (x"c7",x"fe",x"a2",x"49"),
   469 => (x"9f",x"69",x"49",x"ca"),
   470 => (x"e9",x"d5",x"a9",x"02"),
   471 => (x"c0",x"cc",x"87",x"c0"),
   472 => (x"e5",x"ed",x"49",x"d7"),
   473 => (x"cd",x"87",x"c0",x"48"),
   474 => (x"c7",x"fe",x"87",x"73"),
   475 => (x"1e",x"c0",x"e6",x"cb"),
   476 => (x"1e",x"c0",x"e2",x"db"),
   477 => (x"87",x"c1",x"c2",x"d6"),
   478 => (x"1e",x"73",x"49",x"f7"),
   479 => (x"f8",x"87",x"cc",x"86"),
   480 => (x"70",x"98",x"05",x"c0"),
   481 => (x"c5",x"87",x"c0",x"48"),
   482 => (x"c7",x"de",x"87",x"c0"),
   483 => (x"e6",x"e3",x"49",x"d6"),
   484 => (x"e1",x"87",x"c0",x"e8"),
   485 => (x"eb",x"1e",x"c0",x"e1"),
   486 => (x"f6",x"87",x"c8",x"1e"),
   487 => (x"c0",x"e9",x"c3",x"1e"),
   488 => (x"c1",x"c3",x"e8",x"49"),
   489 => (x"fa",x"e2",x"87",x"cc"),
   490 => (x"86",x"70",x"98",x"05"),
   491 => (x"c0",x"c9",x"87",x"c1"),
   492 => (x"ca",x"de",x"48",x"c1"),
   493 => (x"78",x"c0",x"e4",x"87"),
   494 => (x"c8",x"1e",x"c0",x"e9"),
   495 => (x"cc",x"1e",x"c1",x"c3"),
   496 => (x"cc",x"49",x"fa",x"c4"),
   497 => (x"87",x"c8",x"86",x"70"),
   498 => (x"98",x"02",x"c0",x"cf"),
   499 => (x"87",x"c0",x"e7",x"ca"),
   500 => (x"1e",x"c0",x"e0",x"fb"),
   501 => (x"87",x"c4",x"86",x"c0"),
   502 => (x"48",x"c6",x"cd",x"87"),
   503 => (x"c1",x"ca",x"d4",x"97"),
   504 => (x"bf",x"49",x"c1",x"d5"),
   505 => (x"a9",x"05",x"c0",x"cd"),
   506 => (x"87",x"c1",x"ca",x"d5"),
   507 => (x"97",x"bf",x"49",x"c2"),
   508 => (x"ea",x"a9",x"02",x"c0"),
   509 => (x"c5",x"87",x"c0",x"48"),
   510 => (x"c5",x"ee",x"87",x"c1"),
   511 => (x"c2",x"d6",x"97",x"bf"),
   512 => (x"49",x"c3",x"e9",x"a9"),
   513 => (x"02",x"c0",x"d2",x"87"),
   514 => (x"c1",x"c2",x"d6",x"97"),
   515 => (x"bf",x"49",x"c3",x"eb"),
   516 => (x"a9",x"02",x"c0",x"c5"),
   517 => (x"87",x"c0",x"48",x"c5"),
   518 => (x"cf",x"87",x"c1",x"c2"),
   519 => (x"e1",x"97",x"bf",x"49"),
   520 => (x"71",x"99",x"05",x"c0"),
   521 => (x"cc",x"87",x"c1",x"c2"),
   522 => (x"e2",x"97",x"bf",x"49"),
   523 => (x"c2",x"a9",x"02",x"c0"),
   524 => (x"c5",x"87",x"c0",x"48"),
   525 => (x"c4",x"f2",x"87",x"c1"),
   526 => (x"c2",x"e3",x"97",x"bf"),
   527 => (x"48",x"c1",x"ca",x"da"),
   528 => (x"58",x"c1",x"ca",x"d6"),
   529 => (x"bf",x"48",x"c1",x"88"),
   530 => (x"c1",x"ca",x"de",x"58"),
   531 => (x"c1",x"c2",x"e4",x"97"),
   532 => (x"bf",x"49",x"73",x"81"),
   533 => (x"c1",x"c2",x"e5",x"97"),
   534 => (x"bf",x"4a",x"c8",x"32"),
   535 => (x"c1",x"ca",x"ea",x"48"),
   536 => (x"72",x"a1",x"78",x"c1"),
   537 => (x"c2",x"e6",x"97",x"bf"),
   538 => (x"48",x"c1",x"cb",x"c2"),
   539 => (x"58",x"c1",x"ca",x"de"),
   540 => (x"bf",x"02",x"c2",x"e2"),
   541 => (x"87",x"c8",x"1e",x"c0"),
   542 => (x"e7",x"e7",x"1e",x"c1"),
   543 => (x"c3",x"e8",x"49",x"f7"),
   544 => (x"c7",x"87",x"c8",x"86"),
   545 => (x"70",x"98",x"02",x"c0"),
   546 => (x"c5",x"87",x"c0",x"48"),
   547 => (x"c3",x"da",x"87",x"c1"),
   548 => (x"ca",x"d6",x"bf",x"48"),
   549 => (x"c4",x"30",x"c1",x"cb"),
   550 => (x"c6",x"58",x"c1",x"ca"),
   551 => (x"d6",x"bf",x"4a",x"c1"),
   552 => (x"ca",x"fe",x"5a",x"c1"),
   553 => (x"c2",x"fb",x"97",x"bf"),
   554 => (x"49",x"c8",x"31",x"c1"),
   555 => (x"c2",x"fa",x"97",x"bf"),
   556 => (x"4b",x"73",x"a1",x"49"),
   557 => (x"c1",x"c2",x"fc",x"97"),
   558 => (x"bf",x"4b",x"d0",x"33"),
   559 => (x"73",x"a1",x"49",x"c1"),
   560 => (x"c2",x"fd",x"97",x"bf"),
   561 => (x"4b",x"d8",x"33",x"73"),
   562 => (x"a1",x"49",x"c1",x"cb"),
   563 => (x"ca",x"59",x"c1",x"ca"),
   564 => (x"fe",x"bf",x"91",x"c1"),
   565 => (x"ca",x"ea",x"bf",x"81"),
   566 => (x"c1",x"ca",x"f2",x"59"),
   567 => (x"c1",x"c3",x"c3",x"97"),
   568 => (x"bf",x"4b",x"c8",x"33"),
   569 => (x"c1",x"c3",x"c2",x"97"),
   570 => (x"bf",x"4c",x"74",x"a3"),
   571 => (x"4b",x"c1",x"c3",x"c4"),
   572 => (x"97",x"bf",x"4c",x"d0"),
   573 => (x"34",x"74",x"a3",x"4b"),
   574 => (x"c1",x"c3",x"c5",x"97"),
   575 => (x"bf",x"4c",x"cf",x"9c"),
   576 => (x"d8",x"34",x"74",x"a3"),
   577 => (x"4b",x"c1",x"ca",x"f6"),
   578 => (x"5b",x"c2",x"8b",x"73"),
   579 => (x"92",x"c1",x"ca",x"f6"),
   580 => (x"48",x"72",x"a1",x"78"),
   581 => (x"c1",x"d0",x"87",x"c1"),
   582 => (x"c2",x"e8",x"97",x"bf"),
   583 => (x"49",x"c8",x"31",x"c1"),
   584 => (x"c2",x"e7",x"97",x"bf"),
   585 => (x"4a",x"72",x"a1",x"49"),
   586 => (x"c1",x"cb",x"c6",x"59"),
   587 => (x"c5",x"31",x"c7",x"ff"),
   588 => (x"81",x"c9",x"29",x"c1"),
   589 => (x"ca",x"fe",x"59",x"c1"),
   590 => (x"c2",x"ed",x"97",x"bf"),
   591 => (x"4a",x"c8",x"32",x"c1"),
   592 => (x"c2",x"ec",x"97",x"bf"),
   593 => (x"4b",x"73",x"a2",x"4a"),
   594 => (x"c1",x"cb",x"ca",x"5a"),
   595 => (x"c1",x"ca",x"fe",x"bf"),
   596 => (x"92",x"c1",x"ca",x"ea"),
   597 => (x"bf",x"82",x"c1",x"ca"),
   598 => (x"fa",x"5a",x"c1",x"ca"),
   599 => (x"f2",x"48",x"c0",x"78"),
   600 => (x"c1",x"ca",x"ee",x"48"),
   601 => (x"72",x"a1",x"78",x"c1"),
   602 => (x"48",x"26",x"f4",x"d8"),
   603 => (x"87",x"4e",x"6f",x"20"),
   604 => (x"70",x"61",x"72",x"74"),
   605 => (x"69",x"74",x"69",x"6f"),
   606 => (x"6e",x"20",x"73",x"69"),
   607 => (x"67",x"6e",x"61",x"74"),
   608 => (x"75",x"72",x"65",x"20"),
   609 => (x"66",x"6f",x"75",x"6e"),
   610 => (x"64",x"0a",x"00",x"52"),
   611 => (x"65",x"61",x"64",x"69"),
   612 => (x"6e",x"67",x"20",x"62"),
   613 => (x"6f",x"6f",x"74",x"20"),
   614 => (x"73",x"65",x"63",x"74"),
   615 => (x"6f",x"72",x"20",x"25"),
   616 => (x"64",x"0a",x"00",x"52"),
   617 => (x"65",x"61",x"64",x"20"),
   618 => (x"62",x"6f",x"6f",x"74"),
   619 => (x"20",x"73",x"65",x"63"),
   620 => (x"74",x"6f",x"72",x"20"),
   621 => (x"66",x"72",x"6f",x"6d"),
   622 => (x"20",x"66",x"69",x"72"),
   623 => (x"73",x"74",x"20",x"70"),
   624 => (x"61",x"72",x"74",x"69"),
   625 => (x"74",x"69",x"6f",x"6e"),
   626 => (x"0a",x"00",x"55",x"6e"),
   627 => (x"73",x"75",x"70",x"70"),
   628 => (x"6f",x"72",x"74",x"65"),
   629 => (x"64",x"20",x"70",x"61"),
   630 => (x"72",x"74",x"69",x"74"),
   631 => (x"69",x"6f",x"6e",x"20"),
   632 => (x"74",x"79",x"70",x"65"),
   633 => (x"21",x"0d",x"00",x"46"),
   634 => (x"41",x"54",x"33",x"32"),
   635 => (x"20",x"20",x"20",x"00"),
   636 => (x"52",x"65",x"61",x"64"),
   637 => (x"69",x"6e",x"67",x"20"),
   638 => (x"4d",x"42",x"52",x"0a"),
   639 => (x"00",x"46",x"41",x"54"),
   640 => (x"31",x"36",x"20",x"20"),
   641 => (x"20",x"00",x"46",x"41"),
   642 => (x"54",x"33",x"32",x"20"),
   643 => (x"20",x"20",x"00",x"46"),
   644 => (x"41",x"54",x"31",x"32"),
   645 => (x"20",x"20",x"20",x"00"),
   646 => (x"50",x"61",x"72",x"74"),
   647 => (x"69",x"74",x"69",x"6f"),
   648 => (x"6e",x"63",x"6f",x"75"),
   649 => (x"6e",x"74",x"20",x"25"),
   650 => (x"64",x"0a",x"00",x"48"),
   651 => (x"75",x"6e",x"74",x"69"),
   652 => (x"6e",x"67",x"20",x"66"),
   653 => (x"6f",x"72",x"20",x"66"),
   654 => (x"69",x"6c",x"65",x"73"),
   655 => (x"79",x"73",x"74",x"65"),
   656 => (x"6d",x"0a",x"00",x"46"),
   657 => (x"41",x"54",x"33",x"32"),
   658 => (x"20",x"20",x"20",x"00"),
   659 => (x"46",x"41",x"54",x"31"),
   660 => (x"36",x"20",x"20",x"20"),
   661 => (x"00",x"52",x"65",x"61"),
   662 => (x"64",x"69",x"6e",x"67"),
   663 => (x"20",x"64",x"69",x"72"),
   664 => (x"65",x"63",x"74",x"6f"),
   665 => (x"72",x"79",x"20",x"73"),
   666 => (x"65",x"63",x"74",x"6f"),
   667 => (x"72",x"20",x"25",x"64"),
   668 => (x"0a",x"00",x"66",x"69"),
   669 => (x"6c",x"65",x"20",x"22"),
   670 => (x"25",x"73",x"22",x"20"),
   671 => (x"66",x"6f",x"75",x"6e"),
   672 => (x"64",x"0d",x"00",x"47"),
   673 => (x"65",x"74",x"46",x"41"),
   674 => (x"54",x"4c",x"69",x"6e"),
   675 => (x"6b",x"20",x"72",x"65"),
   676 => (x"74",x"75",x"72",x"6e"),
   677 => (x"65",x"64",x"20",x"25"),
   678 => (x"64",x"0a",x"00",x"43"),
   679 => (x"61",x"6e",x"27",x"74"),
   680 => (x"20",x"6f",x"70",x"65"),
   681 => (x"6e",x"20",x"25",x"73"),
   682 => (x"0a",x"00",x"0e",x"5e"),
   683 => (x"5b",x"5c",x"5d",x"0e"),
   684 => (x"71",x"4a",x"c1",x"ca"),
   685 => (x"de",x"bf",x"02",x"cc"),
   686 => (x"87",x"72",x"4b",x"c7"),
   687 => (x"b7",x"2b",x"72",x"4c"),
   688 => (x"c1",x"ff",x"9c",x"ca"),
   689 => (x"87",x"72",x"4b",x"c8"),
   690 => (x"b7",x"2b",x"72",x"4c"),
   691 => (x"c3",x"ff",x"9c",x"c1"),
   692 => (x"cb",x"ce",x"bf",x"ab"),
   693 => (x"02",x"de",x"87",x"c1"),
   694 => (x"c2",x"d6",x"1e",x"c1"),
   695 => (x"ca",x"ea",x"bf",x"49"),
   696 => (x"73",x"81",x"ea",x"d1"),
   697 => (x"87",x"c4",x"86",x"70"),
   698 => (x"98",x"05",x"c5",x"87"),
   699 => (x"c0",x"48",x"c0",x"f6"),
   700 => (x"87",x"c1",x"cb",x"d2"),
   701 => (x"5b",x"c1",x"ca",x"de"),
   702 => (x"bf",x"02",x"d9",x"87"),
   703 => (x"74",x"4a",x"c4",x"92"),
   704 => (x"c1",x"c2",x"d6",x"82"),
   705 => (x"6a",x"49",x"eb",x"ec"),
   706 => (x"87",x"70",x"49",x"71"),
   707 => (x"4d",x"cf",x"ff",x"ff"),
   708 => (x"ff",x"ff",x"9d",x"d0"),
   709 => (x"87",x"74",x"4a",x"c2"),
   710 => (x"92",x"c1",x"c2",x"d6"),
   711 => (x"82",x"9f",x"6a",x"49"),
   712 => (x"ec",x"cc",x"87",x"70"),
   713 => (x"4d",x"75",x"48",x"ed"),
   714 => (x"d9",x"87",x"0e",x"5e"),
   715 => (x"5b",x"5c",x"5d",x"0e"),
   716 => (x"f4",x"86",x"71",x"4c"),
   717 => (x"c0",x"4b",x"c1",x"cb"),
   718 => (x"ce",x"48",x"ff",x"78"),
   719 => (x"c1",x"ca",x"f2",x"bf"),
   720 => (x"4d",x"c1",x"ca",x"f6"),
   721 => (x"bf",x"7e",x"c1",x"ca"),
   722 => (x"de",x"bf",x"02",x"c9"),
   723 => (x"87",x"c1",x"ca",x"d6"),
   724 => (x"bf",x"4a",x"c4",x"32"),
   725 => (x"c7",x"87",x"c1",x"ca"),
   726 => (x"fa",x"bf",x"4a",x"c4"),
   727 => (x"32",x"c8",x"a6",x"5a"),
   728 => (x"c8",x"a6",x"48",x"c0"),
   729 => (x"78",x"c4",x"66",x"48"),
   730 => (x"c0",x"a8",x"06",x"c3"),
   731 => (x"cf",x"87",x"c8",x"66"),
   732 => (x"49",x"cf",x"99",x"05"),
   733 => (x"c0",x"e3",x"87",x"6e"),
   734 => (x"1e",x"c0",x"e9",x"d5"),
   735 => (x"1e",x"d2",x"d0",x"87"),
   736 => (x"c1",x"c2",x"d6",x"1e"),
   737 => (x"cc",x"66",x"49",x"48"),
   738 => (x"c1",x"80",x"d0",x"a6"),
   739 => (x"58",x"71",x"49",x"e7"),
   740 => (x"e4",x"87",x"cc",x"86"),
   741 => (x"c1",x"c2",x"d6",x"4b"),
   742 => (x"c3",x"87",x"c0",x"e0"),
   743 => (x"83",x"97",x"6b",x"49"),
   744 => (x"71",x"99",x"02",x"c2"),
   745 => (x"c5",x"87",x"97",x"6b"),
   746 => (x"49",x"c3",x"e5",x"a9"),
   747 => (x"02",x"c1",x"fb",x"87"),
   748 => (x"cb",x"a3",x"49",x"97"),
   749 => (x"69",x"49",x"d8",x"99"),
   750 => (x"05",x"c1",x"ef",x"87"),
   751 => (x"cb",x"1e",x"c0",x"e0"),
   752 => (x"66",x"1e",x"73",x"49"),
   753 => (x"ea",x"c2",x"87",x"c8"),
   754 => (x"86",x"70",x"98",x"05"),
   755 => (x"c1",x"dc",x"87",x"dc"),
   756 => (x"a3",x"4a",x"6a",x"49"),
   757 => (x"e8",x"de",x"87",x"70"),
   758 => (x"4a",x"c4",x"a4",x"49"),
   759 => (x"72",x"79",x"da",x"a3"),
   760 => (x"4a",x"9f",x"6a",x"49"),
   761 => (x"e9",x"c8",x"87",x"c4"),
   762 => (x"a6",x"58",x"c1",x"ca"),
   763 => (x"de",x"bf",x"02",x"d8"),
   764 => (x"87",x"d4",x"a3",x"4a"),
   765 => (x"9f",x"6a",x"49",x"e8"),
   766 => (x"f5",x"87",x"70",x"49"),
   767 => (x"c0",x"ff",x"ff",x"99"),
   768 => (x"71",x"48",x"d0",x"30"),
   769 => (x"c8",x"a6",x"58",x"c5"),
   770 => (x"87",x"c4",x"a6",x"48"),
   771 => (x"c0",x"78",x"c4",x"66"),
   772 => (x"4a",x"6e",x"82",x"c8"),
   773 => (x"a4",x"49",x"72",x"79"),
   774 => (x"c0",x"7c",x"dc",x"66"),
   775 => (x"1e",x"c0",x"e9",x"f2"),
   776 => (x"1e",x"cf",x"ec",x"87"),
   777 => (x"c8",x"86",x"c1",x"48"),
   778 => (x"c1",x"d0",x"87",x"c8"),
   779 => (x"66",x"48",x"c1",x"80"),
   780 => (x"cc",x"a6",x"58",x"c8"),
   781 => (x"66",x"48",x"c4",x"66"),
   782 => (x"a8",x"04",x"fc",x"f1"),
   783 => (x"87",x"c1",x"ca",x"de"),
   784 => (x"bf",x"02",x"c0",x"f4"),
   785 => (x"87",x"75",x"49",x"f9"),
   786 => (x"e0",x"87",x"70",x"4d"),
   787 => (x"75",x"1e",x"c0",x"ea"),
   788 => (x"c3",x"1e",x"ce",x"fb"),
   789 => (x"87",x"c8",x"86",x"75"),
   790 => (x"49",x"cf",x"ff",x"ff"),
   791 => (x"ff",x"f8",x"99",x"a9"),
   792 => (x"02",x"d6",x"87",x"75"),
   793 => (x"49",x"c2",x"89",x"c1"),
   794 => (x"ca",x"d6",x"bf",x"91"),
   795 => (x"c1",x"ca",x"ee",x"bf"),
   796 => (x"48",x"71",x"80",x"c4"),
   797 => (x"a6",x"58",x"fb",x"e7"),
   798 => (x"87",x"c0",x"48",x"f4"),
   799 => (x"8e",x"e8",x"c3",x"87"),
   800 => (x"0e",x"5e",x"5b",x"5c"),
   801 => (x"5d",x"0e",x"1e",x"71"),
   802 => (x"4b",x"73",x"1e",x"c1"),
   803 => (x"cb",x"d2",x"49",x"fa"),
   804 => (x"d8",x"87",x"c4",x"86"),
   805 => (x"70",x"98",x"02",x"c1"),
   806 => (x"f7",x"87",x"c1",x"cb"),
   807 => (x"d6",x"bf",x"49",x"c7"),
   808 => (x"ff",x"81",x"c9",x"29"),
   809 => (x"c4",x"a6",x"59",x"c0"),
   810 => (x"4d",x"4c",x"6e",x"48"),
   811 => (x"c0",x"b7",x"a8",x"06"),
   812 => (x"c1",x"ed",x"87",x"c1"),
   813 => (x"ca",x"ee",x"bf",x"49"),
   814 => (x"c1",x"cb",x"da",x"bf"),
   815 => (x"4a",x"c2",x"8a",x"c1"),
   816 => (x"ca",x"d6",x"bf",x"92"),
   817 => (x"72",x"a1",x"49",x"c1"),
   818 => (x"ca",x"da",x"bf",x"4a"),
   819 => (x"74",x"9a",x"72",x"a1"),
   820 => (x"49",x"d4",x"66",x"1e"),
   821 => (x"71",x"49",x"e2",x"dd"),
   822 => (x"87",x"c4",x"86",x"70"),
   823 => (x"98",x"05",x"c5",x"87"),
   824 => (x"c0",x"48",x"c1",x"c0"),
   825 => (x"87",x"c1",x"84",x"c1"),
   826 => (x"ca",x"da",x"bf",x"49"),
   827 => (x"74",x"99",x"05",x"cc"),
   828 => (x"87",x"c1",x"cb",x"da"),
   829 => (x"bf",x"49",x"f6",x"f1"),
   830 => (x"87",x"c1",x"cb",x"de"),
   831 => (x"58",x"d4",x"66",x"48"),
   832 => (x"c8",x"c0",x"80",x"d8"),
   833 => (x"a6",x"58",x"c1",x"85"),
   834 => (x"6e",x"b7",x"ad",x"04"),
   835 => (x"fe",x"e4",x"87",x"cf"),
   836 => (x"87",x"73",x"1e",x"c0"),
   837 => (x"ea",x"db",x"1e",x"cb"),
   838 => (x"f6",x"87",x"c8",x"86"),
   839 => (x"c0",x"48",x"c5",x"87"),
   840 => (x"c1",x"cb",x"d6",x"bf"),
   841 => (x"48",x"26",x"e5",x"da"),
   842 => (x"87",x"1e",x"f3",x"09"),
   843 => (x"97",x"79",x"09",x"71"),
   844 => (x"48",x"26",x"4f",x"0e"),
   845 => (x"5e",x"5b",x"5c",x"0e"),
   846 => (x"71",x"4b",x"c0",x"4c"),
   847 => (x"13",x"4a",x"72",x"9a"),
   848 => (x"02",x"cd",x"87",x"72"),
   849 => (x"49",x"e2",x"87",x"c1"),
   850 => (x"84",x"13",x"4a",x"72"),
   851 => (x"9a",x"05",x"f3",x"87"),
   852 => (x"74",x"48",x"c2",x"87"),
   853 => (x"26",x"4d",x"26",x"4c"),
   854 => (x"26",x"4b",x"26",x"4f"),
   855 => (x"0e",x"5e",x"5b",x"5c"),
   856 => (x"5d",x"0e",x"fc",x"86"),
   857 => (x"71",x"4a",x"c0",x"e0"),
   858 => (x"66",x"4c",x"c1",x"cb"),
   859 => (x"de",x"4b",x"c0",x"7e"),
   860 => (x"72",x"9a",x"05",x"ce"),
   861 => (x"87",x"c1",x"cb",x"df"),
   862 => (x"4b",x"c1",x"cb",x"de"),
   863 => (x"48",x"c0",x"f0",x"50"),
   864 => (x"c1",x"d2",x"87",x"72"),
   865 => (x"9a",x"02",x"c0",x"e9"),
   866 => (x"87",x"d4",x"66",x"4d"),
   867 => (x"72",x"1e",x"72",x"49"),
   868 => (x"75",x"4a",x"ca",x"cf"),
   869 => (x"87",x"26",x"4a",x"c0"),
   870 => (x"f8",x"c6",x"81",x"11"),
   871 => (x"53",x"71",x"1e",x"72"),
   872 => (x"49",x"75",x"4a",x"c9"),
   873 => (x"fe",x"87",x"70",x"4a"),
   874 => (x"26",x"49",x"c1",x"8c"),
   875 => (x"72",x"9a",x"05",x"ff"),
   876 => (x"da",x"87",x"c0",x"b7"),
   877 => (x"ac",x"06",x"dd",x"87"),
   878 => (x"c0",x"e4",x"66",x"02"),
   879 => (x"c5",x"87",x"c0",x"f0"),
   880 => (x"4a",x"c3",x"87",x"c0"),
   881 => (x"e0",x"4a",x"73",x"0a"),
   882 => (x"97",x"7a",x"0a",x"c1"),
   883 => (x"83",x"8c",x"c0",x"b7"),
   884 => (x"ac",x"01",x"ff",x"e3"),
   885 => (x"87",x"c1",x"cb",x"de"),
   886 => (x"ab",x"02",x"de",x"87"),
   887 => (x"d8",x"66",x"4c",x"dc"),
   888 => (x"66",x"1e",x"c1",x"8b"),
   889 => (x"97",x"6b",x"49",x"74"),
   890 => (x"0f",x"c4",x"86",x"6e"),
   891 => (x"48",x"c1",x"80",x"c4"),
   892 => (x"a6",x"58",x"c1",x"cb"),
   893 => (x"de",x"ab",x"05",x"ff"),
   894 => (x"e5",x"87",x"6e",x"48"),
   895 => (x"fc",x"8e",x"26",x"4d"),
   896 => (x"26",x"4c",x"26",x"4b"),
   897 => (x"26",x"4f",x"30",x"31"),
   898 => (x"32",x"33",x"34",x"35"),
   899 => (x"36",x"37",x"38",x"39"),
   900 => (x"41",x"42",x"43",x"44"),
   901 => (x"45",x"46",x"00",x"0e"),
   902 => (x"5e",x"5b",x"5c",x"5d"),
   903 => (x"0e",x"71",x"4b",x"ff"),
   904 => (x"4d",x"13",x"4c",x"74"),
   905 => (x"9c",x"02",x"d8",x"87"),
   906 => (x"c1",x"85",x"d4",x"66"),
   907 => (x"1e",x"74",x"49",x"d4"),
   908 => (x"66",x"0f",x"c4",x"86"),
   909 => (x"74",x"a8",x"05",x"c7"),
   910 => (x"87",x"13",x"4c",x"74"),
   911 => (x"9c",x"05",x"e8",x"87"),
   912 => (x"75",x"48",x"26",x"4d"),
   913 => (x"26",x"4c",x"26",x"4b"),
   914 => (x"26",x"4f",x"0e",x"5e"),
   915 => (x"5b",x"5c",x"5d",x"0e"),
   916 => (x"e8",x"86",x"c4",x"a6"),
   917 => (x"59",x"c0",x"e8",x"66"),
   918 => (x"4d",x"c0",x"4c",x"c8"),
   919 => (x"a6",x"48",x"c0",x"78"),
   920 => (x"6e",x"97",x"bf",x"4b"),
   921 => (x"6e",x"48",x"c1",x"80"),
   922 => (x"c4",x"a6",x"58",x"73"),
   923 => (x"9b",x"02",x"c6",x"d3"),
   924 => (x"87",x"c8",x"66",x"02"),
   925 => (x"c5",x"db",x"87",x"cc"),
   926 => (x"a6",x"48",x"c0",x"78"),
   927 => (x"fc",x"80",x"c0",x"78"),
   928 => (x"73",x"4a",x"c0",x"e0"),
   929 => (x"8a",x"02",x"c3",x"c6"),
   930 => (x"87",x"c3",x"8a",x"02"),
   931 => (x"c3",x"c0",x"87",x"c2"),
   932 => (x"8a",x"02",x"c2",x"e8"),
   933 => (x"87",x"c2",x"8a",x"02"),
   934 => (x"c2",x"f4",x"87",x"c4"),
   935 => (x"8a",x"02",x"c2",x"ee"),
   936 => (x"87",x"c2",x"8a",x"02"),
   937 => (x"c2",x"e8",x"87",x"c3"),
   938 => (x"8a",x"02",x"c2",x"ea"),
   939 => (x"87",x"d4",x"8a",x"02"),
   940 => (x"c0",x"f6",x"87",x"d4"),
   941 => (x"8a",x"02",x"c1",x"c0"),
   942 => (x"87",x"ca",x"8a",x"02"),
   943 => (x"c0",x"f2",x"87",x"c1"),
   944 => (x"8a",x"02",x"c1",x"e1"),
   945 => (x"87",x"c1",x"8a",x"02"),
   946 => (x"df",x"87",x"c8",x"8a"),
   947 => (x"02",x"c1",x"ce",x"87"),
   948 => (x"c4",x"8a",x"02",x"c0"),
   949 => (x"e3",x"87",x"c3",x"8a"),
   950 => (x"02",x"c0",x"e5",x"87"),
   951 => (x"c2",x"8a",x"02",x"c8"),
   952 => (x"87",x"c3",x"8a",x"02"),
   953 => (x"d3",x"87",x"c1",x"fa"),
   954 => (x"87",x"cc",x"a6",x"48"),
   955 => (x"ca",x"78",x"c2",x"d2"),
   956 => (x"87",x"cc",x"a6",x"48"),
   957 => (x"c2",x"78",x"c2",x"ca"),
   958 => (x"87",x"cc",x"a6",x"48"),
   959 => (x"d0",x"78",x"c2",x"c2"),
   960 => (x"87",x"c0",x"f0",x"66"),
   961 => (x"1e",x"c0",x"f0",x"66"),
   962 => (x"1e",x"c4",x"85",x"75"),
   963 => (x"4a",x"c4",x"8a",x"6a"),
   964 => (x"49",x"fc",x"c3",x"87"),
   965 => (x"c8",x"86",x"70",x"49"),
   966 => (x"71",x"a4",x"4c",x"c1"),
   967 => (x"e5",x"87",x"c8",x"a6"),
   968 => (x"48",x"c1",x"78",x"c1"),
   969 => (x"dd",x"87",x"c0",x"f0"),
   970 => (x"66",x"1e",x"c4",x"85"),
   971 => (x"75",x"4a",x"c4",x"8a"),
   972 => (x"6a",x"49",x"c0",x"f0"),
   973 => (x"66",x"0f",x"c4",x"86"),
   974 => (x"c1",x"84",x"c1",x"c6"),
   975 => (x"87",x"c0",x"f0",x"66"),
   976 => (x"1e",x"c0",x"e5",x"49"),
   977 => (x"c0",x"f0",x"66",x"0f"),
   978 => (x"c4",x"86",x"c1",x"84"),
   979 => (x"c0",x"f4",x"87",x"c8"),
   980 => (x"a6",x"48",x"c1",x"78"),
   981 => (x"c0",x"ec",x"87",x"d0"),
   982 => (x"a6",x"48",x"c1",x"78"),
   983 => (x"f8",x"80",x"c1",x"78"),
   984 => (x"c0",x"e0",x"87",x"c0"),
   985 => (x"f0",x"ab",x"06",x"da"),
   986 => (x"87",x"c0",x"f9",x"ab"),
   987 => (x"03",x"d4",x"87",x"d4"),
   988 => (x"66",x"49",x"ca",x"91"),
   989 => (x"73",x"4a",x"c0",x"f0"),
   990 => (x"8a",x"d4",x"a6",x"48"),
   991 => (x"72",x"a1",x"78",x"f4"),
   992 => (x"80",x"c1",x"78",x"cc"),
   993 => (x"66",x"02",x"c1",x"ea"),
   994 => (x"87",x"c4",x"85",x"75"),
   995 => (x"49",x"c4",x"89",x"a6"),
   996 => (x"48",x"69",x"78",x"c1"),
   997 => (x"e4",x"ab",x"05",x"d8"),
   998 => (x"87",x"c4",x"66",x"48"),
   999 => (x"c0",x"b7",x"a8",x"03"),
  1000 => (x"cf",x"87",x"c0",x"ed"),
  1001 => (x"49",x"f6",x"c1",x"87"),
  1002 => (x"c4",x"66",x"48",x"c0"),
  1003 => (x"08",x"88",x"c8",x"a6"),
  1004 => (x"58",x"d0",x"66",x"1e"),
  1005 => (x"d8",x"66",x"1e",x"c0"),
  1006 => (x"f8",x"66",x"1e",x"c0"),
  1007 => (x"f8",x"66",x"1e",x"dc"),
  1008 => (x"66",x"1e",x"d8",x"66"),
  1009 => (x"49",x"f6",x"d4",x"87"),
  1010 => (x"d4",x"86",x"70",x"49"),
  1011 => (x"71",x"a4",x"4c",x"c0"),
  1012 => (x"e1",x"87",x"c0",x"e5"),
  1013 => (x"ab",x"05",x"cf",x"87"),
  1014 => (x"d0",x"a6",x"48",x"c0"),
  1015 => (x"78",x"c4",x"80",x"c0"),
  1016 => (x"78",x"f4",x"80",x"c1"),
  1017 => (x"78",x"cc",x"87",x"c0"),
  1018 => (x"f0",x"66",x"1e",x"73"),
  1019 => (x"49",x"c0",x"f0",x"66"),
  1020 => (x"0f",x"c4",x"86",x"6e"),
  1021 => (x"97",x"bf",x"4b",x"6e"),
  1022 => (x"48",x"c1",x"80",x"c4"),
  1023 => (x"a6",x"58",x"73",x"9b"),
  1024 => (x"05",x"f9",x"ed",x"87"),
  1025 => (x"74",x"48",x"e8",x"8e"),
  1026 => (x"26",x"4d",x"26",x"4c"),
  1027 => (x"26",x"4b",x"26",x"4f"),
  1028 => (x"1e",x"c0",x"1e",x"c0"),
  1029 => (x"f4",x"e9",x"1e",x"d0"),
  1030 => (x"a6",x"1e",x"d0",x"66"),
  1031 => (x"49",x"f8",x"ea",x"87"),
  1032 => (x"f4",x"8e",x"26",x"4f"),
  1033 => (x"1e",x"73",x"1e",x"72"),
  1034 => (x"9a",x"02",x"c0",x"e7"),
  1035 => (x"87",x"c0",x"48",x"c1"),
  1036 => (x"4b",x"72",x"a9",x"06"),
  1037 => (x"d1",x"87",x"72",x"82"),
  1038 => (x"06",x"c9",x"87",x"73"),
  1039 => (x"83",x"72",x"a9",x"01"),
  1040 => (x"f4",x"87",x"c3",x"87"),
  1041 => (x"c1",x"b2",x"3a",x"72"),
  1042 => (x"a9",x"03",x"89",x"73"),
  1043 => (x"80",x"07",x"c1",x"2a"),
  1044 => (x"2b",x"05",x"f3",x"87"),
  1045 => (x"26",x"4b",x"26",x"4f"),
  1046 => (x"1e",x"75",x"1e",x"c4"),
  1047 => (x"4d",x"71",x"b7",x"a1"),
  1048 => (x"04",x"ff",x"b9",x"c1"),
  1049 => (x"81",x"c3",x"bd",x"07"),
  1050 => (x"72",x"b7",x"a2",x"04"),
  1051 => (x"ff",x"ba",x"c1",x"82"),
  1052 => (x"c1",x"bd",x"07",x"fe"),
  1053 => (x"ee",x"87",x"c1",x"2d"),
  1054 => (x"04",x"ff",x"b8",x"c1"),
  1055 => (x"80",x"07",x"2d",x"04"),
  1056 => (x"ff",x"b9",x"c1",x"81"),
  1057 => (x"07",x"26",x"4d",x"26"),
  1058 => (x"4f",x"26",x"4d",x"26"),
	others => (others => x"00")
);

-- Xilinx XST attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "no_rw_check";

-- Altera Quartus attributes
attribute ramstyle: string;
attribute ramstyle of ram: signal is "no_rw_check";

signal q_local : word_t;

begin
    
	process(clk,q_local)
	begin

		q(31 downto 24)<=q_local(0);
		q(23 downto 16)<=q_local(1);
		q(15 downto 8)<=q_local(2);
		q(7 downto 0)<=q_local(3);

		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel(3) = '1') then
					ram(to_integer(unsigned(addr)))(3) <= d(7 downto 0);
				end if;
				if bytesel(2) = '1' then
					ram(to_integer(unsigned(addr)))(2) <= d(15 downto 8);
				end if;
				if bytesel(1) = '1' then
					ram(to_integer(unsigned(addr)))(1) <= d(23 downto 16);
				end if;
				if bytesel(0) = '1' then
					ram(to_integer(unsigned(addr)))(0) <= d(31 downto 24);
				end if;
			end if;
			q_local <= ram(to_integer(unsigned(addr)));
		end if;
	end process;

end arch;

