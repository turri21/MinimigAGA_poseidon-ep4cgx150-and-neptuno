library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM-2 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111";
	-- Second port
	addr2 : in std_logic_vector(maxAddrBitBRAM-2 downto 0) := (others=>'0');
	q2 : out std_logic_vector(31 downto 0);
	d2 : in std_logic_vector(31 downto 0) := X"00000000";
	we2 : in std_logic := '0';
	bytesel2 : in std_logic_vector(3 downto 0) := "1111"	
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
type ram_type is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

signal ram : ram_type :=
(
     0 => (x"01",x"da",x"87",x"04"),
     1 => (x"dd",x"87",x"0e",x"58"),
     2 => (x"5e",x"59",x"5a",x"0e"),
     3 => (x"27",x"00",x"00",x"00"),
     4 => (x"29",x"0f",x"26",x"4a"),
     5 => (x"26",x"49",x"26",x"48"),
     6 => (x"ff",x"80",x"26",x"08"),
     7 => (x"4f",x"27",x"00",x"00"),
     8 => (x"00",x"2d",x"4f",x"27"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"4f",x"4f",x"00",x"fd"),
    11 => (x"87",x"c1",x"cd",x"d4"),
    12 => (x"4e",x"c9",x"c0",x"86"),
    13 => (x"c1",x"cd",x"d4",x"49"),
    14 => (x"c1",x"c3",x"f0",x"48"),
    15 => (x"89",x"d0",x"89",x"03"),
    16 => (x"c0",x"40",x"40",x"40"),
    17 => (x"40",x"f6",x"87",x"d0"),
    18 => (x"81",x"05",x"c0",x"50"),
    19 => (x"c1",x"89",x"05",x"f9"),
    20 => (x"87",x"c1",x"c3",x"ed"),
    21 => (x"4d",x"c1",x"c3",x"ed"),
    22 => (x"4c",x"74",x"ad",x"02"),
    23 => (x"c4",x"87",x"24",x"0f"),
    24 => (x"f7",x"87",x"c2",x"df"),
    25 => (x"87",x"c1",x"c3",x"ed"),
    26 => (x"4d",x"c1",x"c3",x"ed"),
    27 => (x"4c",x"74",x"ad",x"02"),
    28 => (x"c6",x"87",x"c4",x"8c"),
    29 => (x"6c",x"0f",x"f5",x"87"),
    30 => (x"00",x"fd",x"87",x"0e"),
    31 => (x"5e",x"5b",x"5c",x"0e"),
    32 => (x"c4",x"c0",x"c0",x"c0"),
    33 => (x"4b",x"c9",x"c3",x"4c"),
    34 => (x"c9",x"d5",x"bf",x"4a"),
    35 => (x"49",x"c1",x"8a",x"71"),
    36 => (x"99",x"02",x"cf",x"87"),
    37 => (x"74",x"49",x"c1",x"84"),
    38 => (x"11",x"53",x"72",x"49"),
    39 => (x"c1",x"8a",x"71",x"99"),
    40 => (x"05",x"f1",x"87",x"c2"),
    41 => (x"87",x"26",x"4d",x"26"),
    42 => (x"4c",x"26",x"4b",x"26"),
    43 => (x"4f",x"1e",x"73",x"1e"),
    44 => (x"71",x"4b",x"e7",x"48"),
    45 => (x"c0",x"e0",x"50",x"e3"),
    46 => (x"48",x"c8",x"50",x"e3"),
    47 => (x"48",x"c6",x"50",x"e7"),
    48 => (x"48",x"c0",x"e1",x"50"),
    49 => (x"73",x"4a",x"c8",x"b7"),
    50 => (x"2a",x"c4",x"c0",x"c0"),
    51 => (x"c0",x"49",x"ca",x"81"),
    52 => (x"71",x"0a",x"97",x"7a"),
    53 => (x"73",x"4a",x"c3",x"ff"),
    54 => (x"9a",x"c4",x"c0",x"c0"),
    55 => (x"c0",x"49",x"cb",x"81"),
    56 => (x"71",x"0a",x"97",x"7a"),
    57 => (x"e7",x"48",x"c0",x"e0"),
    58 => (x"50",x"e3",x"48",x"c8"),
    59 => (x"50",x"e3",x"48",x"c0"),
    60 => (x"50",x"e7",x"48",x"c0"),
    61 => (x"e1",x"50",x"fe",x"f0"),
    62 => (x"87",x"1e",x"73",x"1e"),
    63 => (x"c2",x"c0",x"c0",x"4b"),
    64 => (x"0f",x"fe",x"e5",x"87"),
    65 => (x"1e",x"73",x"1e",x"eb"),
    66 => (x"48",x"c3",x"ef",x"50"),
    67 => (x"e7",x"48",x"c0",x"e0"),
    68 => (x"50",x"e3",x"48",x"c8"),
    69 => (x"50",x"e3",x"48",x"c6"),
    70 => (x"50",x"e7",x"48",x"c0"),
    71 => (x"e1",x"50",x"ff",x"c2"),
    72 => (x"48",x"c1",x"9f",x"78"),
    73 => (x"e7",x"48",x"c0",x"e0"),
    74 => (x"50",x"e3",x"48",x"c4"),
    75 => (x"50",x"e3",x"48",x"c2"),
    76 => (x"50",x"e7",x"48",x"c0"),
    77 => (x"e1",x"50",x"e7",x"48"),
    78 => (x"c0",x"e0",x"50",x"e3"),
    79 => (x"48",x"c8",x"50",x"e3"),
    80 => (x"48",x"c7",x"50",x"e7"),
    81 => (x"48",x"c0",x"e1",x"50"),
    82 => (x"fc",x"f0",x"87",x"c0"),
    83 => (x"ff",x"ff",x"49",x"fd"),
    84 => (x"db",x"87",x"c0",x"fc"),
    85 => (x"c0",x"4b",x"c8",x"cf"),
    86 => (x"49",x"c0",x"f1",x"c7"),
    87 => (x"87",x"d0",x"eb",x"87"),
    88 => (x"70",x"98",x"02",x"c1"),
    89 => (x"c3",x"87",x"c0",x"ff"),
    90 => (x"f0",x"4b",x"c7",x"f8"),
    91 => (x"49",x"c0",x"f0",x"f3"),
    92 => (x"87",x"d6",x"d8",x"87"),
    93 => (x"70",x"98",x"02",x"c0"),
    94 => (x"e6",x"87",x"c3",x"f0"),
    95 => (x"4b",x"c2",x"c0",x"c0"),
    96 => (x"1e",x"c6",x"fb",x"49"),
    97 => (x"c0",x"ed",x"eb",x"87"),
    98 => (x"c4",x"86",x"70",x"98"),
    99 => (x"02",x"c8",x"87",x"c3"),
   100 => (x"ff",x"4b",x"fd",x"e4"),
   101 => (x"87",x"d9",x"87",x"c7"),
   102 => (x"c7",x"49",x"c0",x"f0"),
   103 => (x"c6",x"87",x"d0",x"87"),
   104 => (x"c7",x"dc",x"49",x"c0"),
   105 => (x"ef",x"fd",x"87",x"c7"),
   106 => (x"87",x"c8",x"e5",x"49"),
   107 => (x"c0",x"ef",x"f4",x"87"),
   108 => (x"73",x"49",x"fb",x"f8"),
   109 => (x"87",x"fe",x"da",x"87"),
   110 => (x"fb",x"ee",x"87",x"38"),
   111 => (x"33",x"32",x"4f",x"53"),
   112 => (x"44",x"41",x"44",x"42"),
   113 => (x"49",x"4e",x"00",x"43"),
   114 => (x"61",x"6e",x"27",x"74"),
   115 => (x"20",x"6c",x"6f",x"61"),
   116 => (x"64",x"20",x"66",x"69"),
   117 => (x"72",x"6d",x"77",x"61"),
   118 => (x"72",x"65",x"0a",x"00"),
   119 => (x"55",x"6e",x"61",x"62"),
   120 => (x"6c",x"65",x"20",x"74"),
   121 => (x"6f",x"20",x"6c",x"6f"),
   122 => (x"63",x"61",x"74",x"65"),
   123 => (x"20",x"70",x"61",x"72"),
   124 => (x"74",x"69",x"74",x"69"),
   125 => (x"6f",x"6e",x"0a",x"00"),
   126 => (x"48",x"75",x"6e",x"74"),
   127 => (x"69",x"6e",x"67",x"20"),
   128 => (x"66",x"6f",x"72",x"20"),
   129 => (x"70",x"61",x"72",x"74"),
   130 => (x"69",x"74",x"69",x"6f"),
   131 => (x"6e",x"0a",x"00",x"49"),
   132 => (x"6e",x"69",x"74",x"69"),
   133 => (x"61",x"6c",x"69",x"7a"),
   134 => (x"69",x"6e",x"67",x"20"),
   135 => (x"53",x"44",x"20",x"63"),
   136 => (x"61",x"72",x"64",x"0a"),
   137 => (x"00",x"46",x"61",x"69"),
   138 => (x"6c",x"65",x"64",x"20"),
   139 => (x"74",x"6f",x"20",x"69"),
   140 => (x"6e",x"69",x"74",x"69"),
   141 => (x"61",x"6c",x"69",x"7a"),
   142 => (x"65",x"20",x"53",x"44"),
   143 => (x"20",x"63",x"61",x"72"),
   144 => (x"64",x"0a",x"00",x"00"),
   145 => (x"00",x"00",x"00",x"00"),
   146 => (x"00",x"00",x"08",x"33"),
   147 => (x"fc",x"0f",x"ff",x"00"),
   148 => (x"df",x"f1",x"80",x"60"),
   149 => (x"f6",x"00",x"00",x"00"),
   150 => (x"12",x"1e",x"e4",x"86"),
   151 => (x"e3",x"48",x"c3",x"ff"),
   152 => (x"50",x"e3",x"97",x"bf"),
   153 => (x"48",x"c4",x"a6",x"58"),
   154 => (x"70",x"49",x"c3",x"ff"),
   155 => (x"99",x"e3",x"48",x"c3"),
   156 => (x"ff",x"50",x"c8",x"31"),
   157 => (x"e3",x"97",x"bf",x"48"),
   158 => (x"c8",x"a6",x"58",x"c3"),
   159 => (x"ff",x"98",x"cc",x"a6"),
   160 => (x"58",x"70",x"b1",x"e3"),
   161 => (x"48",x"c3",x"ff",x"50"),
   162 => (x"c8",x"31",x"e3",x"97"),
   163 => (x"bf",x"48",x"d0",x"a6"),
   164 => (x"58",x"c3",x"ff",x"98"),
   165 => (x"d4",x"a6",x"58",x"70"),
   166 => (x"b1",x"e3",x"48",x"c3"),
   167 => (x"ff",x"50",x"c8",x"31"),
   168 => (x"e3",x"97",x"bf",x"48"),
   169 => (x"d8",x"a6",x"58",x"c3"),
   170 => (x"ff",x"98",x"dc",x"a6"),
   171 => (x"58",x"70",x"b1",x"71"),
   172 => (x"48",x"e4",x"8e",x"26"),
   173 => (x"4f",x"0e",x"5e",x"5b"),
   174 => (x"5c",x"0e",x"1e",x"71"),
   175 => (x"4a",x"49",x"c3",x"ff"),
   176 => (x"99",x"e3",x"09",x"97"),
   177 => (x"79",x"09",x"c1",x"c3"),
   178 => (x"f0",x"bf",x"05",x"c8"),
   179 => (x"87",x"d0",x"66",x"48"),
   180 => (x"c9",x"30",x"d4",x"a6"),
   181 => (x"58",x"d0",x"66",x"49"),
   182 => (x"d8",x"29",x"c3",x"ff"),
   183 => (x"99",x"e3",x"09",x"97"),
   184 => (x"79",x"09",x"d0",x"66"),
   185 => (x"49",x"d0",x"29",x"c3"),
   186 => (x"ff",x"99",x"e3",x"09"),
   187 => (x"97",x"79",x"09",x"d0"),
   188 => (x"66",x"49",x"c8",x"29"),
   189 => (x"c3",x"ff",x"99",x"e3"),
   190 => (x"09",x"97",x"79",x"09"),
   191 => (x"d0",x"66",x"49",x"c3"),
   192 => (x"ff",x"99",x"e3",x"09"),
   193 => (x"97",x"79",x"09",x"72"),
   194 => (x"49",x"d0",x"29",x"c3"),
   195 => (x"ff",x"99",x"e3",x"09"),
   196 => (x"97",x"79",x"09",x"97"),
   197 => (x"bf",x"48",x"c4",x"a6"),
   198 => (x"58",x"70",x"4b",x"c3"),
   199 => (x"ff",x"9b",x"c9",x"f0"),
   200 => (x"ff",x"4c",x"c3",x"ff"),
   201 => (x"ab",x"05",x"dc",x"87"),
   202 => (x"e3",x"48",x"c3",x"ff"),
   203 => (x"50",x"e3",x"97",x"bf"),
   204 => (x"48",x"c4",x"a6",x"58"),
   205 => (x"70",x"4b",x"c3",x"ff"),
   206 => (x"9b",x"c1",x"8c",x"02"),
   207 => (x"c6",x"87",x"c3",x"ff"),
   208 => (x"ab",x"02",x"e4",x"87"),
   209 => (x"73",x"4a",x"c4",x"b7"),
   210 => (x"2a",x"c0",x"f0",x"a2"),
   211 => (x"49",x"c0",x"e9",x"c9"),
   212 => (x"87",x"73",x"4a",x"cf"),
   213 => (x"9a",x"c0",x"f0",x"a2"),
   214 => (x"49",x"c0",x"e8",x"fd"),
   215 => (x"87",x"73",x"48",x"26"),
   216 => (x"c2",x"87",x"26",x"4d"),
   217 => (x"26",x"4c",x"26",x"4b"),
   218 => (x"26",x"4f",x"1e",x"c0"),
   219 => (x"49",x"e3",x"48",x"c3"),
   220 => (x"ff",x"50",x"c1",x"81"),
   221 => (x"c3",x"c8",x"b7",x"a9"),
   222 => (x"04",x"f2",x"87",x"26"),
   223 => (x"4f",x"1e",x"73",x"1e"),
   224 => (x"e8",x"87",x"c4",x"f8"),
   225 => (x"df",x"4b",x"c0",x"1e"),
   226 => (x"c0",x"ff",x"f0",x"c1"),
   227 => (x"f7",x"49",x"fc",x"e4"),
   228 => (x"87",x"c4",x"86",x"c1"),
   229 => (x"a8",x"05",x"c0",x"e8"),
   230 => (x"87",x"e3",x"48",x"c3"),
   231 => (x"ff",x"50",x"c1",x"c0"),
   232 => (x"c0",x"c0",x"c0",x"c0"),
   233 => (x"1e",x"c0",x"e1",x"f0"),
   234 => (x"c1",x"e9",x"49",x"fc"),
   235 => (x"c7",x"87",x"c4",x"86"),
   236 => (x"70",x"98",x"05",x"c9"),
   237 => (x"87",x"e3",x"48",x"c3"),
   238 => (x"ff",x"50",x"c1",x"48"),
   239 => (x"cb",x"87",x"fe",x"e9"),
   240 => (x"87",x"c1",x"8b",x"05"),
   241 => (x"fe",x"ff",x"87",x"c0"),
   242 => (x"48",x"fe",x"da",x"87"),
   243 => (x"43",x"4d",x"44",x"34"),
   244 => (x"31",x"20",x"25",x"64"),
   245 => (x"0a",x"00",x"43",x"4d"),
   246 => (x"44",x"35",x"35",x"20"),
   247 => (x"25",x"64",x"0a",x"00"),
   248 => (x"43",x"4d",x"44",x"34"),
   249 => (x"31",x"20",x"25",x"64"),
   250 => (x"0a",x"00",x"43",x"4d"),
   251 => (x"44",x"35",x"35",x"20"),
   252 => (x"25",x"64",x"0a",x"00"),
   253 => (x"69",x"6e",x"69",x"74"),
   254 => (x"20",x"25",x"64",x"0a"),
   255 => (x"20",x"20",x"00",x"69"),
   256 => (x"6e",x"69",x"74",x"20"),
   257 => (x"25",x"64",x"0a",x"20"),
   258 => (x"20",x"00",x"43",x"6d"),
   259 => (x"64",x"5f",x"69",x"6e"),
   260 => (x"69",x"74",x"0a",x"00"),
   261 => (x"43",x"4d",x"44",x"38"),
   262 => (x"5f",x"34",x"20",x"72"),
   263 => (x"65",x"73",x"70",x"6f"),
   264 => (x"6e",x"73",x"65",x"3a"),
   265 => (x"20",x"25",x"64",x"0a"),
   266 => (x"00",x"43",x"4d",x"44"),
   267 => (x"35",x"38",x"20",x"25"),
   268 => (x"64",x"0a",x"20",x"20"),
   269 => (x"00",x"43",x"4d",x"44"),
   270 => (x"35",x"38",x"5f",x"32"),
   271 => (x"20",x"25",x"64",x"0a"),
   272 => (x"20",x"20",x"00",x"43"),
   273 => (x"4d",x"44",x"35",x"38"),
   274 => (x"20",x"25",x"64",x"0a"),
   275 => (x"20",x"20",x"00",x"53"),
   276 => (x"44",x"48",x"43",x"20"),
   277 => (x"49",x"6e",x"69",x"74"),
   278 => (x"69",x"61",x"6c",x"69"),
   279 => (x"7a",x"61",x"74",x"69"),
   280 => (x"6f",x"6e",x"20",x"65"),
   281 => (x"72",x"72",x"6f",x"72"),
   282 => (x"21",x"0a",x"00",x"63"),
   283 => (x"6d",x"64",x"5f",x"43"),
   284 => (x"4d",x"44",x"38",x"20"),
   285 => (x"72",x"65",x"73",x"70"),
   286 => (x"6f",x"6e",x"73",x"65"),
   287 => (x"3a",x"20",x"25",x"64"),
   288 => (x"0a",x"00",x"52",x"65"),
   289 => (x"61",x"64",x"20",x"63"),
   290 => (x"6f",x"6d",x"6d",x"61"),
   291 => (x"6e",x"64",x"20",x"66"),
   292 => (x"61",x"69",x"6c",x"65"),
   293 => (x"64",x"20",x"61",x"74"),
   294 => (x"20",x"25",x"64",x"20"),
   295 => (x"28",x"25",x"64",x"29"),
   296 => (x"0a",x"00",x"1e",x"73"),
   297 => (x"1e",x"e3",x"48",x"c3"),
   298 => (x"ff",x"50",x"d0",x"ca"),
   299 => (x"49",x"c0",x"e3",x"f3"),
   300 => (x"87",x"d3",x"4b",x"c0"),
   301 => (x"1e",x"c0",x"ff",x"f0"),
   302 => (x"c1",x"c1",x"49",x"f7"),
   303 => (x"f7",x"87",x"c4",x"86"),
   304 => (x"70",x"98",x"05",x"c9"),
   305 => (x"87",x"e3",x"48",x"c3"),
   306 => (x"ff",x"50",x"c1",x"48"),
   307 => (x"cb",x"87",x"fa",x"d9"),
   308 => (x"87",x"c1",x"8b",x"05"),
   309 => (x"ff",x"dc",x"87",x"c0"),
   310 => (x"48",x"fa",x"ca",x"87"),
   311 => (x"1e",x"73",x"1e",x"1e"),
   312 => (x"fa",x"c7",x"87",x"c6"),
   313 => (x"ea",x"1e",x"c0",x"e1"),
   314 => (x"f0",x"c1",x"c8",x"49"),
   315 => (x"f7",x"c6",x"87",x"70"),
   316 => (x"4b",x"1e",x"d1",x"eb"),
   317 => (x"1e",x"c0",x"ed",x"fb"),
   318 => (x"87",x"cc",x"86",x"c1"),
   319 => (x"ab",x"02",x"c8",x"87"),
   320 => (x"fe",x"df",x"87",x"c0"),
   321 => (x"48",x"c1",x"ff",x"87"),
   322 => (x"f5",x"ce",x"87",x"70"),
   323 => (x"49",x"cf",x"ff",x"ff"),
   324 => (x"99",x"c6",x"ea",x"a9"),
   325 => (x"02",x"c8",x"87",x"fe"),
   326 => (x"c8",x"87",x"c0",x"48"),
   327 => (x"c1",x"e8",x"87",x"e3"),
   328 => (x"48",x"c3",x"ff",x"50"),
   329 => (x"c0",x"f1",x"4b",x"f9"),
   330 => (x"d3",x"87",x"70",x"98"),
   331 => (x"02",x"c1",x"c6",x"87"),
   332 => (x"c0",x"1e",x"c0",x"ff"),
   333 => (x"f0",x"c1",x"fa",x"49"),
   334 => (x"f5",x"fa",x"87",x"c4"),
   335 => (x"86",x"70",x"98",x"05"),
   336 => (x"c0",x"f3",x"87",x"e3"),
   337 => (x"48",x"c3",x"ff",x"50"),
   338 => (x"e3",x"97",x"bf",x"48"),
   339 => (x"c4",x"a6",x"58",x"70"),
   340 => (x"49",x"c3",x"ff",x"99"),
   341 => (x"e3",x"48",x"c3",x"ff"),
   342 => (x"50",x"e3",x"48",x"c3"),
   343 => (x"ff",x"50",x"e3",x"48"),
   344 => (x"c3",x"ff",x"50",x"e3"),
   345 => (x"48",x"c3",x"ff",x"50"),
   346 => (x"c1",x"c0",x"99",x"02"),
   347 => (x"c4",x"87",x"c1",x"48"),
   348 => (x"d5",x"87",x"c0",x"48"),
   349 => (x"d1",x"87",x"c2",x"ab"),
   350 => (x"05",x"c4",x"87",x"c0"),
   351 => (x"48",x"c8",x"87",x"c1"),
   352 => (x"8b",x"05",x"fe",x"e2"),
   353 => (x"87",x"c0",x"48",x"26"),
   354 => (x"f7",x"db",x"87",x"1e"),
   355 => (x"73",x"1e",x"c1",x"c3"),
   356 => (x"f0",x"48",x"c1",x"78"),
   357 => (x"eb",x"48",x"c3",x"ef"),
   358 => (x"50",x"c7",x"4b",x"e7"),
   359 => (x"48",x"c3",x"50",x"f7"),
   360 => (x"c8",x"87",x"e7",x"48"),
   361 => (x"c2",x"50",x"e3",x"48"),
   362 => (x"c3",x"ff",x"50",x"c0"),
   363 => (x"1e",x"c0",x"e5",x"d0"),
   364 => (x"c1",x"c0",x"49",x"f3"),
   365 => (x"ff",x"87",x"c4",x"86"),
   366 => (x"c1",x"a8",x"05",x"c1"),
   367 => (x"87",x"4b",x"c2",x"ab"),
   368 => (x"05",x"c5",x"87",x"c0"),
   369 => (x"48",x"c0",x"ef",x"87"),
   370 => (x"c1",x"8b",x"05",x"ff"),
   371 => (x"cd",x"87",x"fc",x"cb"),
   372 => (x"87",x"c1",x"c3",x"f4"),
   373 => (x"58",x"70",x"98",x"05"),
   374 => (x"cd",x"87",x"c1",x"1e"),
   375 => (x"c0",x"ff",x"f0",x"c1"),
   376 => (x"d0",x"49",x"f3",x"d0"),
   377 => (x"87",x"c4",x"86",x"e3"),
   378 => (x"48",x"c3",x"ff",x"50"),
   379 => (x"e7",x"48",x"c3",x"50"),
   380 => (x"e3",x"48",x"c3",x"ff"),
   381 => (x"50",x"c1",x"48",x"f5"),
   382 => (x"ec",x"87",x"0e",x"5e"),
   383 => (x"5b",x"5c",x"5d",x"0e"),
   384 => (x"1e",x"71",x"4a",x"c0"),
   385 => (x"4d",x"e3",x"48",x"c3"),
   386 => (x"ff",x"50",x"e7",x"48"),
   387 => (x"c2",x"50",x"eb",x"48"),
   388 => (x"c7",x"50",x"e3",x"48"),
   389 => (x"c3",x"ff",x"50",x"72"),
   390 => (x"1e",x"c0",x"ff",x"f0"),
   391 => (x"c1",x"d1",x"49",x"f2"),
   392 => (x"d3",x"87",x"c4",x"86"),
   393 => (x"70",x"98",x"05",x"c1"),
   394 => (x"c8",x"87",x"c5",x"ee"),
   395 => (x"cd",x"df",x"4b",x"e3"),
   396 => (x"48",x"c3",x"ff",x"50"),
   397 => (x"e3",x"97",x"bf",x"48"),
   398 => (x"c4",x"a6",x"58",x"70"),
   399 => (x"49",x"c3",x"ff",x"99"),
   400 => (x"c3",x"fe",x"a9",x"05"),
   401 => (x"dd",x"87",x"c0",x"4c"),
   402 => (x"f0",x"ce",x"87",x"d4"),
   403 => (x"66",x"08",x"78",x"d4"),
   404 => (x"66",x"48",x"c4",x"80"),
   405 => (x"d8",x"a6",x"58",x"c1"),
   406 => (x"84",x"c2",x"c0",x"b7"),
   407 => (x"ac",x"04",x"e8",x"87"),
   408 => (x"c1",x"4b",x"4d",x"c1"),
   409 => (x"8b",x"05",x"ff",x"c6"),
   410 => (x"87",x"e3",x"48",x"c3"),
   411 => (x"ff",x"50",x"e7",x"48"),
   412 => (x"c3",x"50",x"75",x"48"),
   413 => (x"26",x"f3",x"ea",x"87"),
   414 => (x"1e",x"73",x"1e",x"71"),
   415 => (x"4b",x"49",x"d8",x"29"),
   416 => (x"c3",x"ff",x"99",x"73"),
   417 => (x"4a",x"c8",x"2a",x"cf"),
   418 => (x"fc",x"c0",x"9a",x"72"),
   419 => (x"b1",x"73",x"4a",x"c8"),
   420 => (x"32",x"c0",x"ff",x"f0"),
   421 => (x"c0",x"c0",x"9a",x"72"),
   422 => (x"b1",x"73",x"4a",x"d8"),
   423 => (x"32",x"ff",x"c0",x"c0"),
   424 => (x"c0",x"c0",x"9a",x"72"),
   425 => (x"b1",x"71",x"48",x"c4"),
   426 => (x"87",x"26",x"4d",x"26"),
   427 => (x"4c",x"26",x"4b",x"26"),
   428 => (x"4f",x"1e",x"73",x"1e"),
   429 => (x"71",x"4b",x"49",x"c8"),
   430 => (x"29",x"c3",x"ff",x"99"),
   431 => (x"73",x"4a",x"c8",x"32"),
   432 => (x"cf",x"fc",x"c0",x"9a"),
   433 => (x"72",x"b1",x"71",x"48"),
   434 => (x"e3",x"87",x"0e",x"5e"),
   435 => (x"5b",x"5c",x"0e",x"71"),
   436 => (x"4b",x"c0",x"4c",x"d0"),
   437 => (x"66",x"48",x"c0",x"b7"),
   438 => (x"a8",x"06",x"c0",x"e3"),
   439 => (x"87",x"13",x"4a",x"cc"),
   440 => (x"66",x"97",x"bf",x"49"),
   441 => (x"cc",x"66",x"48",x"c1"),
   442 => (x"80",x"d0",x"a6",x"58"),
   443 => (x"71",x"b7",x"aa",x"02"),
   444 => (x"c4",x"87",x"c1",x"48"),
   445 => (x"cc",x"87",x"c1",x"84"),
   446 => (x"d0",x"66",x"b7",x"ac"),
   447 => (x"04",x"ff",x"dd",x"87"),
   448 => (x"c0",x"48",x"c2",x"87"),
   449 => (x"26",x"4d",x"26",x"4c"),
   450 => (x"26",x"4b",x"26",x"4f"),
   451 => (x"0e",x"5e",x"5b",x"5c"),
   452 => (x"0e",x"1e",x"c1",x"cc"),
   453 => (x"f2",x"48",x"ff",x"78"),
   454 => (x"c1",x"cc",x"c2",x"48"),
   455 => (x"c0",x"78",x"c0",x"e9"),
   456 => (x"e7",x"49",x"d9",x"ff"),
   457 => (x"87",x"c1",x"c3",x"fa"),
   458 => (x"1e",x"c0",x"49",x"fb"),
   459 => (x"cc",x"87",x"c4",x"86"),
   460 => (x"70",x"98",x"05",x"c5"),
   461 => (x"87",x"c0",x"48",x"ca"),
   462 => (x"e6",x"87",x"c0",x"4b"),
   463 => (x"c1",x"cc",x"ee",x"48"),
   464 => (x"c1",x"78",x"c8",x"1e"),
   465 => (x"c0",x"e9",x"f4",x"1e"),
   466 => (x"c1",x"c4",x"f0",x"49"),
   467 => (x"fd",x"fb",x"87",x"c8"),
   468 => (x"86",x"70",x"98",x"05"),
   469 => (x"c6",x"87",x"c1",x"cc"),
   470 => (x"ee",x"48",x"c0",x"78"),
   471 => (x"c8",x"1e",x"c0",x"e9"),
   472 => (x"fd",x"1e",x"c1",x"c5"),
   473 => (x"cc",x"49",x"fd",x"e1"),
   474 => (x"87",x"c8",x"86",x"70"),
   475 => (x"98",x"05",x"c6",x"87"),
   476 => (x"c1",x"cc",x"ee",x"48"),
   477 => (x"c0",x"78",x"c8",x"1e"),
   478 => (x"c0",x"ea",x"c6",x"1e"),
   479 => (x"c1",x"c5",x"cc",x"49"),
   480 => (x"fd",x"c7",x"87",x"c8"),
   481 => (x"86",x"70",x"98",x"05"),
   482 => (x"c5",x"87",x"c0",x"48"),
   483 => (x"c9",x"d1",x"87",x"c1"),
   484 => (x"cc",x"ee",x"bf",x"1e"),
   485 => (x"c0",x"ea",x"cf",x"1e"),
   486 => (x"c0",x"e3",x"d8",x"87"),
   487 => (x"c8",x"86",x"c1",x"cc"),
   488 => (x"ee",x"bf",x"02",x"c1"),
   489 => (x"ed",x"87",x"c1",x"c3"),
   490 => (x"fa",x"4a",x"48",x"c6"),
   491 => (x"fe",x"a0",x"4c",x"c1"),
   492 => (x"cb",x"c0",x"bf",x"4b"),
   493 => (x"c1",x"cb",x"f8",x"9f"),
   494 => (x"bf",x"49",x"c4",x"a6"),
   495 => (x"5a",x"c5",x"d6",x"ea"),
   496 => (x"a9",x"05",x"c0",x"cc"),
   497 => (x"87",x"c8",x"a4",x"4a"),
   498 => (x"6a",x"49",x"fa",x"eb"),
   499 => (x"87",x"70",x"4b",x"db"),
   500 => (x"87",x"c7",x"fe",x"a2"),
   501 => (x"49",x"9f",x"69",x"49"),
   502 => (x"ca",x"e9",x"d5",x"a9"),
   503 => (x"02",x"c0",x"cc",x"87"),
   504 => (x"c0",x"e7",x"e4",x"49"),
   505 => (x"d6",x"fd",x"87",x"c0"),
   506 => (x"48",x"c7",x"f4",x"87"),
   507 => (x"73",x"1e",x"c0",x"e8"),
   508 => (x"c2",x"1e",x"c0",x"e1"),
   509 => (x"fe",x"87",x"c1",x"c3"),
   510 => (x"fa",x"1e",x"73",x"49"),
   511 => (x"f7",x"fb",x"87",x"cc"),
   512 => (x"86",x"70",x"98",x"05"),
   513 => (x"c0",x"c5",x"87",x"c0"),
   514 => (x"48",x"c7",x"d4",x"87"),
   515 => (x"c0",x"e8",x"da",x"49"),
   516 => (x"d6",x"d1",x"87",x"c0"),
   517 => (x"ea",x"e2",x"1e",x"c0"),
   518 => (x"e1",x"d9",x"87",x"c8"),
   519 => (x"1e",x"c0",x"ea",x"fa"),
   520 => (x"1e",x"c1",x"c5",x"cc"),
   521 => (x"49",x"fa",x"e2",x"87"),
   522 => (x"cc",x"86",x"70",x"98"),
   523 => (x"05",x"c0",x"c9",x"87"),
   524 => (x"c1",x"cc",x"c2",x"48"),
   525 => (x"c1",x"78",x"c0",x"e4"),
   526 => (x"87",x"c8",x"1e",x"c0"),
   527 => (x"eb",x"c3",x"1e",x"c1"),
   528 => (x"c4",x"f0",x"49",x"fa"),
   529 => (x"c4",x"87",x"c8",x"86"),
   530 => (x"70",x"98",x"02",x"c0"),
   531 => (x"cf",x"87",x"c0",x"e9"),
   532 => (x"c1",x"1e",x"c0",x"e0"),
   533 => (x"de",x"87",x"c4",x"86"),
   534 => (x"c0",x"48",x"c6",x"c3"),
   535 => (x"87",x"c1",x"cb",x"f8"),
   536 => (x"97",x"bf",x"49",x"c1"),
   537 => (x"d5",x"a9",x"05",x"c0"),
   538 => (x"cd",x"87",x"c1",x"cb"),
   539 => (x"f9",x"97",x"bf",x"49"),
   540 => (x"c2",x"ea",x"a9",x"02"),
   541 => (x"c0",x"c5",x"87",x"c0"),
   542 => (x"48",x"c5",x"e4",x"87"),
   543 => (x"c1",x"c3",x"fa",x"97"),
   544 => (x"bf",x"49",x"c3",x"e9"),
   545 => (x"a9",x"02",x"c0",x"d2"),
   546 => (x"87",x"c1",x"c3",x"fa"),
   547 => (x"97",x"bf",x"49",x"c3"),
   548 => (x"eb",x"a9",x"02",x"c0"),
   549 => (x"c5",x"87",x"c0",x"48"),
   550 => (x"c5",x"c5",x"87",x"c1"),
   551 => (x"c4",x"c5",x"97",x"bf"),
   552 => (x"49",x"99",x"05",x"c0"),
   553 => (x"cc",x"87",x"c1",x"c4"),
   554 => (x"c6",x"97",x"bf",x"49"),
   555 => (x"c2",x"a9",x"02",x"c0"),
   556 => (x"c5",x"87",x"c0",x"48"),
   557 => (x"c4",x"e9",x"87",x"c1"),
   558 => (x"c4",x"c7",x"97",x"bf"),
   559 => (x"48",x"c1",x"cb",x"fe"),
   560 => (x"58",x"c1",x"88",x"c1"),
   561 => (x"cc",x"c2",x"58",x"c1"),
   562 => (x"c4",x"c8",x"97",x"bf"),
   563 => (x"49",x"73",x"81",x"c1"),
   564 => (x"c4",x"c9",x"97",x"bf"),
   565 => (x"4a",x"c8",x"32",x"c1"),
   566 => (x"cc",x"ce",x"48",x"72"),
   567 => (x"a1",x"78",x"c1",x"c4"),
   568 => (x"ca",x"97",x"bf",x"48"),
   569 => (x"c1",x"cc",x"e6",x"58"),
   570 => (x"c1",x"cc",x"c2",x"bf"),
   571 => (x"02",x"c2",x"e0",x"87"),
   572 => (x"c8",x"1e",x"c0",x"e9"),
   573 => (x"de",x"1e",x"c1",x"c5"),
   574 => (x"cc",x"49",x"f7",x"cd"),
   575 => (x"87",x"c8",x"86",x"70"),
   576 => (x"98",x"02",x"c0",x"c5"),
   577 => (x"87",x"c0",x"48",x"c3"),
   578 => (x"d6",x"87",x"c1",x"cb"),
   579 => (x"fa",x"bf",x"48",x"c4"),
   580 => (x"30",x"c1",x"cc",x"ea"),
   581 => (x"58",x"c1",x"cb",x"fa"),
   582 => (x"bf",x"4a",x"c1",x"cc"),
   583 => (x"e2",x"5a",x"c1",x"c4"),
   584 => (x"df",x"97",x"bf",x"49"),
   585 => (x"c8",x"31",x"c1",x"c4"),
   586 => (x"de",x"97",x"bf",x"4b"),
   587 => (x"a1",x"49",x"c1",x"c4"),
   588 => (x"e0",x"97",x"bf",x"4b"),
   589 => (x"d0",x"33",x"73",x"a1"),
   590 => (x"49",x"c1",x"c4",x"e1"),
   591 => (x"97",x"bf",x"4b",x"d8"),
   592 => (x"33",x"73",x"a1",x"49"),
   593 => (x"c1",x"cc",x"ee",x"59"),
   594 => (x"c1",x"cc",x"e2",x"bf"),
   595 => (x"91",x"c1",x"cc",x"ce"),
   596 => (x"bf",x"81",x"c1",x"cc"),
   597 => (x"d6",x"59",x"c1",x"c4"),
   598 => (x"e7",x"97",x"bf",x"4b"),
   599 => (x"c8",x"33",x"c1",x"c4"),
   600 => (x"e6",x"97",x"bf",x"4c"),
   601 => (x"a3",x"4b",x"c1",x"c4"),
   602 => (x"e8",x"97",x"bf",x"4c"),
   603 => (x"d0",x"34",x"74",x"a3"),
   604 => (x"4b",x"c1",x"c4",x"e9"),
   605 => (x"97",x"bf",x"4c",x"cf"),
   606 => (x"9c",x"d8",x"34",x"74"),
   607 => (x"a3",x"4b",x"c1",x"cc"),
   608 => (x"da",x"5b",x"c2",x"8b"),
   609 => (x"73",x"92",x"c1",x"cc"),
   610 => (x"da",x"48",x"72",x"a1"),
   611 => (x"78",x"c1",x"ce",x"87"),
   612 => (x"c1",x"c4",x"cc",x"97"),
   613 => (x"bf",x"49",x"c8",x"31"),
   614 => (x"c1",x"c4",x"cb",x"97"),
   615 => (x"bf",x"4a",x"a1",x"49"),
   616 => (x"c1",x"cc",x"ea",x"59"),
   617 => (x"c5",x"31",x"c7",x"ff"),
   618 => (x"81",x"c9",x"29",x"c1"),
   619 => (x"cc",x"e2",x"59",x"c1"),
   620 => (x"c4",x"d1",x"97",x"bf"),
   621 => (x"4a",x"c8",x"32",x"c1"),
   622 => (x"c4",x"d0",x"97",x"bf"),
   623 => (x"4b",x"a2",x"4a",x"c1"),
   624 => (x"cc",x"ee",x"5a",x"c1"),
   625 => (x"cc",x"e2",x"bf",x"92"),
   626 => (x"c1",x"cc",x"ce",x"bf"),
   627 => (x"82",x"c1",x"cc",x"de"),
   628 => (x"5a",x"c1",x"cc",x"d6"),
   629 => (x"48",x"c0",x"78",x"c1"),
   630 => (x"cc",x"d2",x"48",x"72"),
   631 => (x"a1",x"78",x"c1",x"48"),
   632 => (x"26",x"f4",x"e2",x"87"),
   633 => (x"4e",x"6f",x"20",x"70"),
   634 => (x"61",x"72",x"74",x"69"),
   635 => (x"74",x"69",x"6f",x"6e"),
   636 => (x"20",x"73",x"69",x"67"),
   637 => (x"6e",x"61",x"74",x"75"),
   638 => (x"72",x"65",x"20",x"66"),
   639 => (x"6f",x"75",x"6e",x"64"),
   640 => (x"0a",x"00",x"52",x"65"),
   641 => (x"61",x"64",x"69",x"6e"),
   642 => (x"67",x"20",x"62",x"6f"),
   643 => (x"6f",x"74",x"20",x"73"),
   644 => (x"65",x"63",x"74",x"6f"),
   645 => (x"72",x"20",x"25",x"64"),
   646 => (x"0a",x"00",x"52",x"65"),
   647 => (x"61",x"64",x"20",x"62"),
   648 => (x"6f",x"6f",x"74",x"20"),
   649 => (x"73",x"65",x"63",x"74"),
   650 => (x"6f",x"72",x"20",x"66"),
   651 => (x"72",x"6f",x"6d",x"20"),
   652 => (x"66",x"69",x"72",x"73"),
   653 => (x"74",x"20",x"70",x"61"),
   654 => (x"72",x"74",x"69",x"74"),
   655 => (x"69",x"6f",x"6e",x"0a"),
   656 => (x"00",x"55",x"6e",x"73"),
   657 => (x"75",x"70",x"70",x"6f"),
   658 => (x"72",x"74",x"65",x"64"),
   659 => (x"20",x"70",x"61",x"72"),
   660 => (x"74",x"69",x"74",x"69"),
   661 => (x"6f",x"6e",x"20",x"74"),
   662 => (x"79",x"70",x"65",x"21"),
   663 => (x"0d",x"00",x"46",x"41"),
   664 => (x"54",x"33",x"32",x"20"),
   665 => (x"20",x"20",x"00",x"52"),
   666 => (x"65",x"61",x"64",x"69"),
   667 => (x"6e",x"67",x"20",x"4d"),
   668 => (x"42",x"52",x"0a",x"00"),
   669 => (x"46",x"41",x"54",x"31"),
   670 => (x"36",x"20",x"20",x"20"),
   671 => (x"00",x"46",x"41",x"54"),
   672 => (x"33",x"32",x"20",x"20"),
   673 => (x"20",x"00",x"46",x"41"),
   674 => (x"54",x"31",x"32",x"20"),
   675 => (x"20",x"20",x"00",x"50"),
   676 => (x"61",x"72",x"74",x"69"),
   677 => (x"74",x"69",x"6f",x"6e"),
   678 => (x"63",x"6f",x"75",x"6e"),
   679 => (x"74",x"20",x"25",x"64"),
   680 => (x"0a",x"00",x"48",x"75"),
   681 => (x"6e",x"74",x"69",x"6e"),
   682 => (x"67",x"20",x"66",x"6f"),
   683 => (x"72",x"20",x"66",x"69"),
   684 => (x"6c",x"65",x"73",x"79"),
   685 => (x"73",x"74",x"65",x"6d"),
   686 => (x"0a",x"00",x"46",x"41"),
   687 => (x"54",x"33",x"32",x"20"),
   688 => (x"20",x"20",x"00",x"46"),
   689 => (x"41",x"54",x"31",x"36"),
   690 => (x"20",x"20",x"20",x"00"),
   691 => (x"52",x"65",x"61",x"64"),
   692 => (x"69",x"6e",x"67",x"20"),
   693 => (x"64",x"69",x"72",x"65"),
   694 => (x"63",x"74",x"6f",x"72"),
   695 => (x"79",x"20",x"73",x"65"),
   696 => (x"63",x"74",x"6f",x"72"),
   697 => (x"20",x"25",x"64",x"0a"),
   698 => (x"00",x"66",x"69",x"6c"),
   699 => (x"65",x"20",x"22",x"25"),
   700 => (x"73",x"22",x"20",x"66"),
   701 => (x"6f",x"75",x"6e",x"64"),
   702 => (x"0d",x"00",x"47",x"65"),
   703 => (x"74",x"46",x"41",x"54"),
   704 => (x"4c",x"69",x"6e",x"6b"),
   705 => (x"20",x"72",x"65",x"74"),
   706 => (x"75",x"72",x"6e",x"65"),
   707 => (x"64",x"20",x"25",x"64"),
   708 => (x"0a",x"00",x"43",x"61"),
   709 => (x"6e",x"27",x"74",x"20"),
   710 => (x"6f",x"70",x"65",x"6e"),
   711 => (x"20",x"25",x"73",x"0a"),
   712 => (x"00",x"0e",x"5e",x"5b"),
   713 => (x"5c",x"5d",x"0e",x"71"),
   714 => (x"4a",x"c1",x"cc",x"c2"),
   715 => (x"bf",x"02",x"cc",x"87"),
   716 => (x"72",x"4b",x"c7",x"b7"),
   717 => (x"2b",x"72",x"4c",x"c1"),
   718 => (x"ff",x"9c",x"ca",x"87"),
   719 => (x"72",x"4b",x"c8",x"b7"),
   720 => (x"2b",x"72",x"4c",x"c3"),
   721 => (x"ff",x"9c",x"c1",x"cc"),
   722 => (x"f2",x"bf",x"ab",x"02"),
   723 => (x"de",x"87",x"c1",x"c3"),
   724 => (x"fa",x"1e",x"c1",x"cc"),
   725 => (x"ce",x"bf",x"49",x"73"),
   726 => (x"81",x"ea",x"de",x"87"),
   727 => (x"c4",x"86",x"70",x"98"),
   728 => (x"05",x"c5",x"87",x"c0"),
   729 => (x"48",x"c0",x"f5",x"87"),
   730 => (x"c1",x"cc",x"f6",x"5b"),
   731 => (x"c1",x"cc",x"c2",x"bf"),
   732 => (x"02",x"d8",x"87",x"74"),
   733 => (x"4a",x"c4",x"92",x"c1"),
   734 => (x"c3",x"fa",x"82",x"6a"),
   735 => (x"49",x"eb",x"f8",x"87"),
   736 => (x"70",x"49",x"4d",x"cf"),
   737 => (x"ff",x"ff",x"ff",x"ff"),
   738 => (x"9d",x"d0",x"87",x"74"),
   739 => (x"4a",x"c2",x"92",x"c1"),
   740 => (x"c3",x"fa",x"82",x"9f"),
   741 => (x"6a",x"49",x"ec",x"d8"),
   742 => (x"87",x"70",x"4d",x"75"),
   743 => (x"48",x"ed",x"e4",x"87"),
   744 => (x"0e",x"5e",x"5b",x"5c"),
   745 => (x"5d",x"0e",x"f4",x"86"),
   746 => (x"71",x"4c",x"c0",x"4b"),
   747 => (x"c1",x"cc",x"f2",x"48"),
   748 => (x"ff",x"78",x"c1",x"cc"),
   749 => (x"d6",x"bf",x"4d",x"c1"),
   750 => (x"cc",x"da",x"bf",x"7e"),
   751 => (x"c1",x"cc",x"c2",x"bf"),
   752 => (x"02",x"c9",x"87",x"c1"),
   753 => (x"cb",x"fa",x"bf",x"4a"),
   754 => (x"c4",x"32",x"c7",x"87"),
   755 => (x"c1",x"cc",x"de",x"bf"),
   756 => (x"4a",x"c4",x"32",x"c8"),
   757 => (x"a6",x"5a",x"c8",x"a6"),
   758 => (x"48",x"c0",x"78",x"c4"),
   759 => (x"66",x"48",x"c0",x"a8"),
   760 => (x"06",x"c3",x"cd",x"87"),
   761 => (x"c8",x"66",x"49",x"cf"),
   762 => (x"99",x"05",x"c0",x"e2"),
   763 => (x"87",x"6e",x"1e",x"c0"),
   764 => (x"eb",x"cc",x"1e",x"d1"),
   765 => (x"fe",x"87",x"c1",x"c3"),
   766 => (x"fa",x"1e",x"cc",x"66"),
   767 => (x"49",x"48",x"c1",x"80"),
   768 => (x"d0",x"a6",x"58",x"71"),
   769 => (x"e7",x"f3",x"87",x"cc"),
   770 => (x"86",x"c1",x"c3",x"fa"),
   771 => (x"4b",x"c3",x"87",x"c0"),
   772 => (x"e0",x"83",x"97",x"6b"),
   773 => (x"49",x"99",x"02",x"c2"),
   774 => (x"c5",x"87",x"97",x"6b"),
   775 => (x"49",x"c3",x"e5",x"a9"),
   776 => (x"02",x"c1",x"fb",x"87"),
   777 => (x"cb",x"a3",x"49",x"97"),
   778 => (x"69",x"49",x"d8",x"99"),
   779 => (x"05",x"c1",x"ef",x"87"),
   780 => (x"cb",x"1e",x"c0",x"e0"),
   781 => (x"66",x"1e",x"73",x"49"),
   782 => (x"ea",x"cf",x"87",x"c8"),
   783 => (x"86",x"70",x"98",x"05"),
   784 => (x"c1",x"dc",x"87",x"dc"),
   785 => (x"a3",x"4a",x"6a",x"49"),
   786 => (x"e8",x"ed",x"87",x"70"),
   787 => (x"4a",x"c4",x"a4",x"49"),
   788 => (x"72",x"79",x"da",x"a3"),
   789 => (x"4a",x"9f",x"6a",x"49"),
   790 => (x"e9",x"d6",x"87",x"c4"),
   791 => (x"a6",x"58",x"c1",x"cc"),
   792 => (x"c2",x"bf",x"02",x"d8"),
   793 => (x"87",x"d4",x"a3",x"4a"),
   794 => (x"9f",x"6a",x"49",x"e9"),
   795 => (x"c3",x"87",x"70",x"49"),
   796 => (x"c0",x"ff",x"ff",x"99"),
   797 => (x"71",x"48",x"d0",x"30"),
   798 => (x"c8",x"a6",x"58",x"c5"),
   799 => (x"87",x"c4",x"a6",x"48"),
   800 => (x"c0",x"78",x"c4",x"66"),
   801 => (x"4a",x"6e",x"82",x"c8"),
   802 => (x"a4",x"49",x"72",x"79"),
   803 => (x"c0",x"7c",x"dc",x"66"),
   804 => (x"1e",x"c0",x"eb",x"e9"),
   805 => (x"1e",x"cf",x"dc",x"87"),
   806 => (x"c8",x"86",x"c1",x"48"),
   807 => (x"c1",x"cf",x"87",x"c8"),
   808 => (x"66",x"48",x"c1",x"80"),
   809 => (x"cc",x"a6",x"58",x"c8"),
   810 => (x"66",x"48",x"c4",x"66"),
   811 => (x"a8",x"04",x"fc",x"f3"),
   812 => (x"87",x"c1",x"cc",x"c2"),
   813 => (x"bf",x"02",x"c0",x"f3"),
   814 => (x"87",x"75",x"49",x"f9"),
   815 => (x"e3",x"87",x"70",x"4d"),
   816 => (x"1e",x"c0",x"eb",x"fa"),
   817 => (x"1e",x"ce",x"ec",x"87"),
   818 => (x"c8",x"86",x"75",x"49"),
   819 => (x"cf",x"ff",x"ff",x"ff"),
   820 => (x"f8",x"99",x"a9",x"02"),
   821 => (x"d6",x"87",x"75",x"49"),
   822 => (x"c2",x"89",x"c1",x"cb"),
   823 => (x"fa",x"bf",x"91",x"c1"),
   824 => (x"cc",x"d2",x"bf",x"48"),
   825 => (x"71",x"80",x"c4",x"a6"),
   826 => (x"58",x"fb",x"ea",x"87"),
   827 => (x"c0",x"48",x"f4",x"8e"),
   828 => (x"e8",x"d1",x"87",x"0e"),
   829 => (x"5e",x"5b",x"5c",x"5d"),
   830 => (x"0e",x"1e",x"71",x"4b"),
   831 => (x"1e",x"c1",x"cc",x"f6"),
   832 => (x"49",x"fa",x"dc",x"87"),
   833 => (x"c4",x"86",x"70",x"98"),
   834 => (x"02",x"c1",x"f6",x"87"),
   835 => (x"c1",x"cc",x"fa",x"bf"),
   836 => (x"49",x"c7",x"ff",x"81"),
   837 => (x"c9",x"29",x"c4",x"a6"),
   838 => (x"59",x"c0",x"4d",x"4c"),
   839 => (x"6e",x"48",x"c0",x"b7"),
   840 => (x"a8",x"06",x"c1",x"ec"),
   841 => (x"87",x"c1",x"cc",x"d2"),
   842 => (x"bf",x"49",x"c1",x"cc"),
   843 => (x"fe",x"bf",x"4a",x"c2"),
   844 => (x"8a",x"c1",x"cb",x"fa"),
   845 => (x"bf",x"92",x"72",x"a1"),
   846 => (x"49",x"c1",x"cb",x"fe"),
   847 => (x"bf",x"4a",x"74",x"9a"),
   848 => (x"72",x"a1",x"49",x"d4"),
   849 => (x"66",x"1e",x"71",x"e2"),
   850 => (x"f0",x"87",x"c4",x"86"),
   851 => (x"70",x"98",x"05",x"c5"),
   852 => (x"87",x"c0",x"48",x"c1"),
   853 => (x"c0",x"87",x"c1",x"84"),
   854 => (x"c1",x"cb",x"fe",x"bf"),
   855 => (x"49",x"74",x"99",x"05"),
   856 => (x"cc",x"87",x"c1",x"cc"),
   857 => (x"fe",x"bf",x"49",x"f6"),
   858 => (x"f7",x"87",x"c1",x"cd"),
   859 => (x"c2",x"58",x"d4",x"66"),
   860 => (x"48",x"c8",x"c0",x"80"),
   861 => (x"d8",x"a6",x"58",x"c1"),
   862 => (x"85",x"6e",x"b7",x"ad"),
   863 => (x"04",x"fe",x"e5",x"87"),
   864 => (x"cf",x"87",x"73",x"1e"),
   865 => (x"c0",x"ec",x"d2",x"1e"),
   866 => (x"cb",x"e9",x"87",x"c8"),
   867 => (x"86",x"c0",x"48",x"c5"),
   868 => (x"87",x"c1",x"cc",x"fa"),
   869 => (x"bf",x"48",x"26",x"e5"),
   870 => (x"ea",x"87",x"1e",x"f3"),
   871 => (x"09",x"97",x"79",x"09"),
   872 => (x"71",x"48",x"26",x"4f"),
   873 => (x"0e",x"5e",x"5b",x"5c"),
   874 => (x"0e",x"71",x"4b",x"c0"),
   875 => (x"4c",x"13",x"4a",x"9a"),
   876 => (x"02",x"cc",x"87",x"72"),
   877 => (x"49",x"e3",x"87",x"c1"),
   878 => (x"84",x"13",x"4a",x"9a"),
   879 => (x"05",x"f4",x"87",x"74"),
   880 => (x"48",x"c2",x"87",x"26"),
   881 => (x"4d",x"26",x"4c",x"26"),
   882 => (x"4b",x"26",x"4f",x"0e"),
   883 => (x"5e",x"5b",x"5c",x"5d"),
   884 => (x"0e",x"fc",x"86",x"71"),
   885 => (x"4a",x"c0",x"e0",x"66"),
   886 => (x"4c",x"c1",x"cd",x"c2"),
   887 => (x"4b",x"c0",x"7e",x"72"),
   888 => (x"9a",x"05",x"ce",x"87"),
   889 => (x"c1",x"cd",x"c3",x"4b"),
   890 => (x"c1",x"cd",x"c2",x"48"),
   891 => (x"c0",x"f0",x"50",x"c1"),
   892 => (x"ce",x"87",x"72",x"9a"),
   893 => (x"02",x"c0",x"e5",x"87"),
   894 => (x"d4",x"66",x"4d",x"72"),
   895 => (x"1e",x"72",x"49",x"75"),
   896 => (x"4a",x"ca",x"c4",x"87"),
   897 => (x"26",x"4a",x"c0",x"f9"),
   898 => (x"f1",x"81",x"11",x"53"),
   899 => (x"72",x"49",x"75",x"4a"),
   900 => (x"c9",x"f5",x"87",x"70"),
   901 => (x"4a",x"c1",x"8c",x"72"),
   902 => (x"9a",x"05",x"ff",x"de"),
   903 => (x"87",x"c0",x"b7",x"ac"),
   904 => (x"06",x"dd",x"87",x"c0"),
   905 => (x"e4",x"66",x"02",x"c5"),
   906 => (x"87",x"c0",x"f0",x"4a"),
   907 => (x"c3",x"87",x"c0",x"e0"),
   908 => (x"4a",x"73",x"0a",x"97"),
   909 => (x"7a",x"0a",x"c1",x"83"),
   910 => (x"8c",x"c0",x"b7",x"ac"),
   911 => (x"01",x"ff",x"e3",x"87"),
   912 => (x"c1",x"cd",x"c2",x"ab"),
   913 => (x"02",x"de",x"87",x"d8"),
   914 => (x"66",x"4c",x"dc",x"66"),
   915 => (x"1e",x"c1",x"8b",x"97"),
   916 => (x"6b",x"49",x"74",x"0f"),
   917 => (x"c4",x"86",x"6e",x"48"),
   918 => (x"c1",x"80",x"c4",x"a6"),
   919 => (x"58",x"c1",x"cd",x"c2"),
   920 => (x"ab",x"05",x"ff",x"e5"),
   921 => (x"87",x"6e",x"48",x"fc"),
   922 => (x"8e",x"26",x"4d",x"26"),
   923 => (x"4c",x"26",x"4b",x"26"),
   924 => (x"4f",x"30",x"31",x"32"),
   925 => (x"33",x"34",x"35",x"36"),
   926 => (x"37",x"38",x"39",x"41"),
   927 => (x"42",x"43",x"44",x"45"),
   928 => (x"46",x"00",x"0e",x"5e"),
   929 => (x"5b",x"5c",x"5d",x"0e"),
   930 => (x"71",x"4b",x"ff",x"4d"),
   931 => (x"13",x"4c",x"9c",x"02"),
   932 => (x"d7",x"87",x"c1",x"85"),
   933 => (x"d4",x"66",x"1e",x"74"),
   934 => (x"49",x"d4",x"66",x"0f"),
   935 => (x"c4",x"86",x"74",x"a8"),
   936 => (x"05",x"c6",x"87",x"13"),
   937 => (x"4c",x"9c",x"05",x"e9"),
   938 => (x"87",x"75",x"48",x"26"),
   939 => (x"4d",x"26",x"4c",x"26"),
   940 => (x"4b",x"26",x"4f",x"0e"),
   941 => (x"5e",x"5b",x"5c",x"5d"),
   942 => (x"0e",x"e8",x"86",x"c4"),
   943 => (x"a6",x"59",x"c0",x"e8"),
   944 => (x"66",x"4d",x"c0",x"4c"),
   945 => (x"c8",x"a6",x"48",x"c0"),
   946 => (x"78",x"6e",x"97",x"bf"),
   947 => (x"4b",x"6e",x"48",x"c1"),
   948 => (x"80",x"c4",x"a6",x"58"),
   949 => (x"73",x"9b",x"02",x"c6"),
   950 => (x"ce",x"87",x"c8",x"66"),
   951 => (x"02",x"c5",x"d6",x"87"),
   952 => (x"cc",x"a6",x"48",x"c0"),
   953 => (x"78",x"fc",x"80",x"c0"),
   954 => (x"78",x"73",x"4a",x"c0"),
   955 => (x"e0",x"8a",x"02",x"c3"),
   956 => (x"c2",x"87",x"c3",x"8a"),
   957 => (x"02",x"c2",x"fc",x"87"),
   958 => (x"c2",x"8a",x"02",x"c2"),
   959 => (x"e4",x"87",x"8a",x"02"),
   960 => (x"c2",x"f1",x"87",x"c4"),
   961 => (x"8a",x"02",x"c2",x"eb"),
   962 => (x"87",x"c2",x"8a",x"02"),
   963 => (x"c2",x"e5",x"87",x"c3"),
   964 => (x"8a",x"02",x"c2",x"e7"),
   965 => (x"87",x"d4",x"8a",x"02"),
   966 => (x"c0",x"f4",x"87",x"8a"),
   967 => (x"02",x"c0",x"ff",x"87"),
   968 => (x"ca",x"8a",x"02",x"c0"),
   969 => (x"f1",x"87",x"c1",x"8a"),
   970 => (x"02",x"c1",x"df",x"87"),
   971 => (x"8a",x"02",x"df",x"87"),
   972 => (x"c8",x"8a",x"02",x"c1"),
   973 => (x"cd",x"87",x"c4",x"8a"),
   974 => (x"02",x"c0",x"e3",x"87"),
   975 => (x"c3",x"8a",x"02",x"c0"),
   976 => (x"e5",x"87",x"c2",x"8a"),
   977 => (x"02",x"c8",x"87",x"c3"),
   978 => (x"8a",x"02",x"d3",x"87"),
   979 => (x"c1",x"f9",x"87",x"cc"),
   980 => (x"a6",x"48",x"ca",x"78"),
   981 => (x"c2",x"d1",x"87",x"cc"),
   982 => (x"a6",x"48",x"c2",x"78"),
   983 => (x"c2",x"c9",x"87",x"cc"),
   984 => (x"a6",x"48",x"d0",x"78"),
   985 => (x"c2",x"c1",x"87",x"c0"),
   986 => (x"f0",x"66",x"1e",x"c0"),
   987 => (x"f0",x"66",x"1e",x"c4"),
   988 => (x"85",x"75",x"4a",x"c4"),
   989 => (x"8a",x"6a",x"49",x"fc"),
   990 => (x"c8",x"87",x"c8",x"86"),
   991 => (x"70",x"49",x"a4",x"4c"),
   992 => (x"c1",x"e5",x"87",x"c8"),
   993 => (x"a6",x"48",x"c1",x"78"),
   994 => (x"c1",x"dd",x"87",x"c0"),
   995 => (x"f0",x"66",x"1e",x"c4"),
   996 => (x"85",x"75",x"4a",x"c4"),
   997 => (x"8a",x"6a",x"49",x"c0"),
   998 => (x"f0",x"66",x"0f",x"c4"),
   999 => (x"86",x"c1",x"84",x"c1"),
  1000 => (x"c6",x"87",x"c0",x"f0"),
  1001 => (x"66",x"1e",x"c0",x"e5"),
  1002 => (x"49",x"c0",x"f0",x"66"),
  1003 => (x"0f",x"c4",x"86",x"c1"),
  1004 => (x"84",x"c0",x"f4",x"87"),
  1005 => (x"c8",x"a6",x"48",x"c1"),
  1006 => (x"78",x"c0",x"ec",x"87"),
  1007 => (x"d0",x"a6",x"48",x"c1"),
  1008 => (x"78",x"f8",x"80",x"c1"),
  1009 => (x"78",x"c0",x"e0",x"87"),
  1010 => (x"c0",x"f0",x"ab",x"06"),
  1011 => (x"da",x"87",x"c0",x"f9"),
  1012 => (x"ab",x"03",x"d4",x"87"),
  1013 => (x"d4",x"66",x"49",x"ca"),
  1014 => (x"91",x"73",x"4a",x"c0"),
  1015 => (x"f0",x"8a",x"d4",x"a6"),
  1016 => (x"48",x"72",x"a1",x"78"),
  1017 => (x"f4",x"80",x"c1",x"78"),
  1018 => (x"cc",x"66",x"02",x"c1"),
  1019 => (x"e9",x"87",x"c4",x"85"),
  1020 => (x"75",x"49",x"c4",x"89"),
  1021 => (x"a6",x"48",x"69",x"78"),
  1022 => (x"c1",x"e4",x"ab",x"05"),
  1023 => (x"d8",x"87",x"c4",x"66"),
  1024 => (x"48",x"c0",x"b7",x"a8"),
  1025 => (x"03",x"cf",x"87",x"c0"),
  1026 => (x"ed",x"49",x"f6",x"cd"),
  1027 => (x"87",x"c4",x"66",x"48"),
  1028 => (x"c0",x"08",x"88",x"c8"),
  1029 => (x"a6",x"58",x"d0",x"66"),
  1030 => (x"1e",x"d8",x"66",x"1e"),
  1031 => (x"c0",x"f8",x"66",x"1e"),
  1032 => (x"c0",x"f8",x"66",x"1e"),
  1033 => (x"dc",x"66",x"1e",x"d8"),
  1034 => (x"66",x"49",x"f6",x"de"),
  1035 => (x"87",x"d4",x"86",x"70"),
  1036 => (x"49",x"a4",x"4c",x"c0"),
  1037 => (x"e1",x"87",x"c0",x"e5"),
  1038 => (x"ab",x"05",x"cf",x"87"),
  1039 => (x"d0",x"a6",x"48",x"c0"),
  1040 => (x"78",x"c4",x"80",x"c0"),
  1041 => (x"78",x"f4",x"80",x"c1"),
  1042 => (x"78",x"cc",x"87",x"c0"),
  1043 => (x"f0",x"66",x"1e",x"73"),
  1044 => (x"49",x"c0",x"f0",x"66"),
  1045 => (x"0f",x"c4",x"86",x"6e"),
  1046 => (x"97",x"bf",x"4b",x"6e"),
  1047 => (x"48",x"c1",x"80",x"c4"),
  1048 => (x"a6",x"58",x"73",x"9b"),
  1049 => (x"05",x"f9",x"f2",x"87"),
  1050 => (x"74",x"48",x"e8",x"8e"),
  1051 => (x"26",x"4d",x"26",x"4c"),
  1052 => (x"26",x"4b",x"26",x"4f"),
  1053 => (x"1e",x"c0",x"1e",x"c0"),
  1054 => (x"f6",x"da",x"1e",x"d0"),
  1055 => (x"a6",x"1e",x"d0",x"66"),
  1056 => (x"49",x"f8",x"ef",x"87"),
  1057 => (x"f4",x"8e",x"26",x"4f"),
  1058 => (x"1e",x"73",x"1e",x"72"),
  1059 => (x"9a",x"02",x"c0",x"e7"),
  1060 => (x"87",x"c0",x"48",x"c1"),
  1061 => (x"4b",x"72",x"a9",x"06"),
  1062 => (x"d1",x"87",x"72",x"82"),
  1063 => (x"06",x"c9",x"87",x"73"),
  1064 => (x"83",x"72",x"a9",x"01"),
  1065 => (x"f4",x"87",x"c3",x"87"),
  1066 => (x"c1",x"b2",x"3a",x"72"),
  1067 => (x"a9",x"03",x"89",x"73"),
  1068 => (x"80",x"07",x"c1",x"2a"),
  1069 => (x"2b",x"05",x"f3",x"87"),
  1070 => (x"26",x"4b",x"26",x"4f"),
  1071 => (x"1e",x"75",x"1e",x"c4"),
  1072 => (x"4d",x"71",x"b7",x"a1"),
  1073 => (x"04",x"ff",x"b9",x"c1"),
  1074 => (x"81",x"c3",x"bd",x"07"),
  1075 => (x"72",x"b7",x"a2",x"04"),
  1076 => (x"ff",x"ba",x"c1",x"82"),
  1077 => (x"c1",x"bd",x"07",x"fe"),
  1078 => (x"ee",x"87",x"c1",x"2d"),
  1079 => (x"04",x"ff",x"b8",x"c1"),
  1080 => (x"80",x"07",x"2d",x"04"),
  1081 => (x"ff",x"b9",x"c1",x"81"),
  1082 => (x"07",x"26",x"4d",x"26"),
  1083 => (x"4f",x"26",x"4d",x"26"),
	others => (others => x"00")
);

-- Xilinx XST attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "no_rw_check";

-- Altera Quartus attributes
attribute ramstyle: string;
attribute ramstyle of ram: signal is "no_rw_check";

signal q_local : word_t;
signal q2_local : word_t;

begin
    
	process(clk,q_local)
	begin

		q(31 downto 24)<=q_local(0);
		q(23 downto 16)<=q_local(1);
		q(15 downto 8)<=q_local(2);
		q(7 downto 0)<=q_local(3);

		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel(3) = '1') then
					ram(to_integer(unsigned(addr)))(3) <= d(7 downto 0);
				end if;
				if bytesel(2) = '1' then
					ram(to_integer(unsigned(addr)))(2) <= d(15 downto 8);
				end if;
				if bytesel(1) = '1' then
					ram(to_integer(unsigned(addr)))(1) <= d(23 downto 16);
				end if;
				if bytesel(0) = '1' then
					ram(to_integer(unsigned(addr)))(0) <= d(31 downto 24);
				end if;
			end if;
			q_local <= ram(to_integer(unsigned(addr)));
		end if;
	end process;

	-- Second port
	
	process(clk,q2_local)
	begin

		q2(31 downto 24)<=q2_local(0);
		q2(23 downto 16)<=q2_local(1);
		q2(15 downto 8)<=q2_local(2);
		q2(7 downto 0)<=q2_local(3);

		if(rising_edge(clk)) then 
			if(we2 = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel2(3) = '1') then
					ram(to_integer(unsigned(addr2)))(3) <= d2(7 downto 0);
				end if;
				if bytesel2(2) = '1' then
					ram(to_integer(unsigned(addr2)))(2) <= d2(15 downto 8);
				end if;
				if bytesel2(1) = '1' then
					ram(to_integer(unsigned(addr2)))(1) <= d2(23 downto 16);
				end if;
				if bytesel2(0) = '1' then
					ram(to_integer(unsigned(addr2)))(0) <= d2(31 downto 24);
				end if;
			end if;
			q2_local <= ram(to_integer(unsigned(addr2)));
		end if;
	end process;

end arch;

