library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"01",
     1 => x"da",
     2 => x"87",
     3 => x"04",
     4 => x"dd",
     5 => x"87",
     6 => x"0e",
     7 => x"58",
     8 => x"5e",
     9 => x"59",
    10 => x"5a",
    11 => x"0e",
    12 => x"27",
    13 => x"00",
    14 => x"00",
    15 => x"00",
    16 => x"2c",
    17 => x"0f",
    18 => x"26",
    19 => x"4a",
    20 => x"26",
    21 => x"49",
    22 => x"26",
    23 => x"48",
    24 => x"ff",
    25 => x"80",
    26 => x"26",
    27 => x"08",
    28 => x"4f",
    29 => x"27",
    30 => x"00",
    31 => x"00",
    32 => x"00",
    33 => x"2d",
    34 => x"4f",
    35 => x"27",
    36 => x"00",
    37 => x"00",
    38 => x"00",
    39 => x"29",
    40 => x"4f",
    41 => x"00",
    42 => x"fd",
    43 => x"87",
    44 => x"4f",
    45 => x"c1",
    46 => x"d2",
    47 => x"cc",
    48 => x"4e",
    49 => x"c9",
    50 => x"c0",
    51 => x"86",
    52 => x"c1",
    53 => x"d2",
    54 => x"cc",
    55 => x"49",
    56 => x"c1",
    57 => x"c8",
    58 => x"c8",
    59 => x"48",
    60 => x"89",
    61 => x"d0",
    62 => x"89",
    63 => x"03",
    64 => x"c0",
    65 => x"40",
    66 => x"40",
    67 => x"40",
    68 => x"40",
    69 => x"f6",
    70 => x"87",
    71 => x"d0",
    72 => x"81",
    73 => x"05",
    74 => x"c0",
    75 => x"50",
    76 => x"c1",
    77 => x"89",
    78 => x"05",
    79 => x"f9",
    80 => x"87",
    81 => x"c1",
    82 => x"c8",
    83 => x"c6",
    84 => x"4d",
    85 => x"c1",
    86 => x"c8",
    87 => x"c6",
    88 => x"4c",
    89 => x"74",
    90 => x"ad",
    91 => x"02",
    92 => x"c4",
    93 => x"87",
    94 => x"24",
    95 => x"0f",
    96 => x"f7",
    97 => x"87",
    98 => x"c1",
    99 => x"e6",
   100 => x"87",
   101 => x"c1",
   102 => x"c8",
   103 => x"c6",
   104 => x"4d",
   105 => x"c1",
   106 => x"c8",
   107 => x"c6",
   108 => x"4c",
   109 => x"74",
   110 => x"ad",
   111 => x"02",
   112 => x"c6",
   113 => x"87",
   114 => x"c4",
   115 => x"8c",
   116 => x"6c",
   117 => x"0f",
   118 => x"f5",
   119 => x"87",
   120 => x"00",
   121 => x"fd",
   122 => x"87",
   123 => x"1e",
   124 => x"73",
   125 => x"1e",
   126 => x"c2",
   127 => x"c0",
   128 => x"c0",
   129 => x"4b",
   130 => x"73",
   131 => x"0f",
   132 => x"c4",
   133 => x"87",
   134 => x"26",
   135 => x"4d",
   136 => x"26",
   137 => x"4c",
   138 => x"26",
   139 => x"4b",
   140 => x"26",
   141 => x"4f",
   142 => x"1e",
   143 => x"73",
   144 => x"1e",
   145 => x"c0",
   146 => x"4b",
   147 => x"c8",
   148 => x"66",
   149 => x"4a",
   150 => x"dc",
   151 => x"b7",
   152 => x"2a",
   153 => x"cf",
   154 => x"9a",
   155 => x"c8",
   156 => x"66",
   157 => x"48",
   158 => x"c4",
   159 => x"30",
   160 => x"cc",
   161 => x"a6",
   162 => x"58",
   163 => x"c9",
   164 => x"b7",
   165 => x"aa",
   166 => x"06",
   167 => x"c5",
   168 => x"87",
   169 => x"c0",
   170 => x"f7",
   171 => x"82",
   172 => x"c3",
   173 => x"87",
   174 => x"c0",
   175 => x"f0",
   176 => x"82",
   177 => x"cc",
   178 => x"66",
   179 => x"0a",
   180 => x"97",
   181 => x"7a",
   182 => x"0a",
   183 => x"cc",
   184 => x"66",
   185 => x"48",
   186 => x"c1",
   187 => x"80",
   188 => x"d0",
   189 => x"a6",
   190 => x"58",
   191 => x"c1",
   192 => x"83",
   193 => x"c8",
   194 => x"b7",
   195 => x"ab",
   196 => x"04",
   197 => x"ff",
   198 => x"cb",
   199 => x"87",
   200 => x"fe",
   201 => x"ff",
   202 => x"87",
   203 => x"0e",
   204 => x"5e",
   205 => x"5b",
   206 => x"5c",
   207 => x"5d",
   208 => x"0e",
   209 => x"f0",
   210 => x"86",
   211 => x"c8",
   212 => x"c9",
   213 => x"1e",
   214 => x"c0",
   215 => x"f3",
   216 => x"f2",
   217 => x"87",
   218 => x"c4",
   219 => x"86",
   220 => x"d2",
   221 => x"ce",
   222 => x"87",
   223 => x"70",
   224 => x"98",
   225 => x"02",
   226 => x"c3",
   227 => x"d1",
   228 => x"87",
   229 => x"c7",
   230 => x"f2",
   231 => x"1e",
   232 => x"c0",
   233 => x"f3",
   234 => x"e0",
   235 => x"87",
   236 => x"c4",
   237 => x"86",
   238 => x"d8",
   239 => x"d4",
   240 => x"87",
   241 => x"70",
   242 => x"98",
   243 => x"02",
   244 => x"c2",
   245 => x"f6",
   246 => x"87",
   247 => x"c2",
   248 => x"c0",
   249 => x"c0",
   250 => x"1e",
   251 => x"c7",
   252 => x"ca",
   253 => x"1e",
   254 => x"c0",
   255 => x"f0",
   256 => x"d8",
   257 => x"87",
   258 => x"c8",
   259 => x"86",
   260 => x"70",
   261 => x"4b",
   262 => x"73",
   263 => x"9b",
   264 => x"02",
   265 => x"c2",
   266 => x"ea",
   267 => x"87",
   268 => x"c8",
   269 => x"a6",
   270 => x"48",
   271 => x"c0",
   272 => x"78",
   273 => x"fc",
   274 => x"80",
   275 => x"c2",
   276 => x"c0",
   277 => x"c0",
   278 => x"78",
   279 => x"c0",
   280 => x"4d",
   281 => x"c3",
   282 => x"83",
   283 => x"fc",
   284 => x"9b",
   285 => x"c2",
   286 => x"c0",
   287 => x"c0",
   288 => x"4c",
   289 => x"73",
   290 => x"84",
   291 => x"74",
   292 => x"1e",
   293 => x"c6",
   294 => x"fe",
   295 => x"1e",
   296 => x"c0",
   297 => x"ef",
   298 => x"ee",
   299 => x"87",
   300 => x"c8",
   301 => x"86",
   302 => x"70",
   303 => x"98",
   304 => x"02",
   305 => x"c1",
   306 => x"ef",
   307 => x"87",
   308 => x"c7",
   309 => x"ff",
   310 => x"b7",
   311 => x"ab",
   312 => x"06",
   313 => x"c1",
   314 => x"e7",
   315 => x"87",
   316 => x"c8",
   317 => x"c0",
   318 => x"1e",
   319 => x"c8",
   320 => x"66",
   321 => x"49",
   322 => x"75",
   323 => x"81",
   324 => x"71",
   325 => x"1e",
   326 => x"c0",
   327 => x"f2",
   328 => x"ef",
   329 => x"87",
   330 => x"c8",
   331 => x"86",
   332 => x"70",
   333 => x"49",
   334 => x"d0",
   335 => x"a6",
   336 => x"59",
   337 => x"24",
   338 => x"7e",
   339 => x"c8",
   340 => x"c0",
   341 => x"85",
   342 => x"8b",
   343 => x"cc",
   344 => x"66",
   345 => x"48",
   346 => x"6e",
   347 => x"a8",
   348 => x"02",
   349 => x"c0",
   350 => x"fb",
   351 => x"87",
   352 => x"c8",
   353 => x"66",
   354 => x"48",
   355 => x"c1",
   356 => x"80",
   357 => x"cc",
   358 => x"a6",
   359 => x"58",
   360 => x"c1",
   361 => x"c8",
   362 => x"c8",
   363 => x"1e",
   364 => x"75",
   365 => x"1e",
   366 => x"fc",
   367 => x"dd",
   368 => x"87",
   369 => x"c1",
   370 => x"c8",
   371 => x"d0",
   372 => x"48",
   373 => x"c0",
   374 => x"e0",
   375 => x"50",
   376 => x"c1",
   377 => x"c8",
   378 => x"d1",
   379 => x"1e",
   380 => x"d8",
   381 => x"66",
   382 => x"1e",
   383 => x"fc",
   384 => x"cc",
   385 => x"87",
   386 => x"c1",
   387 => x"c8",
   388 => x"d9",
   389 => x"48",
   390 => x"c0",
   391 => x"e0",
   392 => x"50",
   393 => x"c1",
   394 => x"c8",
   395 => x"da",
   396 => x"1e",
   397 => x"d4",
   398 => x"66",
   399 => x"1e",
   400 => x"fb",
   401 => x"fb",
   402 => x"87",
   403 => x"d8",
   404 => x"86",
   405 => x"c1",
   406 => x"c8",
   407 => x"e2",
   408 => x"48",
   409 => x"c0",
   410 => x"50",
   411 => x"c7",
   412 => x"ff",
   413 => x"b7",
   414 => x"ab",
   415 => x"01",
   416 => x"fe",
   417 => x"d9",
   418 => x"87",
   419 => x"c8",
   420 => x"66",
   421 => x"05",
   422 => x"ce",
   423 => x"87",
   424 => x"fb",
   425 => x"d0",
   426 => x"87",
   427 => x"c9",
   428 => x"87",
   429 => x"c7",
   430 => x"d6",
   431 => x"1e",
   432 => x"c0",
   433 => x"f0",
   434 => x"d8",
   435 => x"87",
   436 => x"c4",
   437 => x"86",
   438 => x"ff",
   439 => x"fd",
   440 => x"87",
   441 => x"f0",
   442 => x"8e",
   443 => x"fb",
   444 => x"c8",
   445 => x"87",
   446 => x"43",
   447 => x"48",
   448 => x"45",
   449 => x"43",
   450 => x"4b",
   451 => x"53",
   452 => x"55",
   453 => x"4d",
   454 => x"42",
   455 => x"49",
   456 => x"4e",
   457 => x"00",
   458 => x"38",
   459 => x"33",
   460 => x"32",
   461 => x"4f",
   462 => x"53",
   463 => x"44",
   464 => x"41",
   465 => x"41",
   466 => x"42",
   467 => x"49",
   468 => x"4e",
   469 => x"00",
   470 => x"55",
   471 => x"6e",
   472 => x"61",
   473 => x"62",
   474 => x"6c",
   475 => x"65",
   476 => x"20",
   477 => x"74",
   478 => x"6f",
   479 => x"20",
   480 => x"6c",
   481 => x"6f",
   482 => x"63",
   483 => x"61",
   484 => x"74",
   485 => x"65",
   486 => x"20",
   487 => x"70",
   488 => x"61",
   489 => x"72",
   490 => x"74",
   491 => x"69",
   492 => x"74",
   493 => x"69",
   494 => x"6f",
   495 => x"6e",
   496 => x"0a",
   497 => x"00",
   498 => x"48",
   499 => x"75",
   500 => x"6e",
   501 => x"74",
   502 => x"69",
   503 => x"6e",
   504 => x"67",
   505 => x"20",
   506 => x"66",
   507 => x"6f",
   508 => x"72",
   509 => x"20",
   510 => x"70",
   511 => x"61",
   512 => x"72",
   513 => x"74",
   514 => x"69",
   515 => x"74",
   516 => x"69",
   517 => x"6f",
   518 => x"6e",
   519 => x"0a",
   520 => x"00",
   521 => x"49",
   522 => x"6e",
   523 => x"69",
   524 => x"74",
   525 => x"69",
   526 => x"61",
   527 => x"6c",
   528 => x"69",
   529 => x"7a",
   530 => x"69",
   531 => x"6e",
   532 => x"67",
   533 => x"20",
   534 => x"53",
   535 => x"44",
   536 => x"20",
   537 => x"63",
   538 => x"61",
   539 => x"72",
   540 => x"64",
   541 => x"0a",
   542 => x"00",
   543 => x"1e",
   544 => x"e4",
   545 => x"86",
   546 => x"c0",
   547 => x"f6",
   548 => x"e4",
   549 => x"c0",
   550 => x"c0",
   551 => x"4a",
   552 => x"c3",
   553 => x"ff",
   554 => x"97",
   555 => x"7a",
   556 => x"97",
   557 => x"6a",
   558 => x"48",
   559 => x"c4",
   560 => x"a6",
   561 => x"58",
   562 => x"6e",
   563 => x"49",
   564 => x"c3",
   565 => x"ff",
   566 => x"99",
   567 => x"97",
   568 => x"7a",
   569 => x"c8",
   570 => x"31",
   571 => x"97",
   572 => x"6a",
   573 => x"48",
   574 => x"c8",
   575 => x"a6",
   576 => x"58",
   577 => x"c4",
   578 => x"66",
   579 => x"48",
   580 => x"c3",
   581 => x"ff",
   582 => x"98",
   583 => x"cc",
   584 => x"a6",
   585 => x"58",
   586 => x"c8",
   587 => x"66",
   588 => x"b1",
   589 => x"c3",
   590 => x"ff",
   591 => x"97",
   592 => x"7a",
   593 => x"c8",
   594 => x"31",
   595 => x"97",
   596 => x"6a",
   597 => x"48",
   598 => x"d0",
   599 => x"a6",
   600 => x"58",
   601 => x"cc",
   602 => x"66",
   603 => x"48",
   604 => x"c3",
   605 => x"ff",
   606 => x"98",
   607 => x"d4",
   608 => x"a6",
   609 => x"58",
   610 => x"d0",
   611 => x"66",
   612 => x"b1",
   613 => x"c3",
   614 => x"ff",
   615 => x"97",
   616 => x"7a",
   617 => x"c8",
   618 => x"31",
   619 => x"12",
   620 => x"48",
   621 => x"d8",
   622 => x"a6",
   623 => x"58",
   624 => x"d4",
   625 => x"66",
   626 => x"48",
   627 => x"c3",
   628 => x"ff",
   629 => x"98",
   630 => x"dc",
   631 => x"a6",
   632 => x"58",
   633 => x"d8",
   634 => x"66",
   635 => x"b1",
   636 => x"71",
   637 => x"48",
   638 => x"e4",
   639 => x"8e",
   640 => x"26",
   641 => x"4f",
   642 => x"0e",
   643 => x"5e",
   644 => x"5b",
   645 => x"5c",
   646 => x"0e",
   647 => x"1e",
   648 => x"c0",
   649 => x"f6",
   650 => x"e4",
   651 => x"c0",
   652 => x"c0",
   653 => x"4b",
   654 => x"d0",
   655 => x"66",
   656 => x"49",
   657 => x"c3",
   658 => x"ff",
   659 => x"99",
   660 => x"73",
   661 => x"09",
   662 => x"97",
   663 => x"79",
   664 => x"09",
   665 => x"c1",
   666 => x"c8",
   667 => x"e8",
   668 => x"bf",
   669 => x"05",
   670 => x"c8",
   671 => x"87",
   672 => x"d4",
   673 => x"66",
   674 => x"48",
   675 => x"c9",
   676 => x"30",
   677 => x"d8",
   678 => x"a6",
   679 => x"58",
   680 => x"d4",
   681 => x"66",
   682 => x"49",
   683 => x"d8",
   684 => x"29",
   685 => x"c3",
   686 => x"ff",
   687 => x"99",
   688 => x"73",
   689 => x"09",
   690 => x"97",
   691 => x"79",
   692 => x"09",
   693 => x"d4",
   694 => x"66",
   695 => x"49",
   696 => x"d0",
   697 => x"29",
   698 => x"c3",
   699 => x"ff",
   700 => x"99",
   701 => x"73",
   702 => x"09",
   703 => x"97",
   704 => x"79",
   705 => x"09",
   706 => x"d4",
   707 => x"66",
   708 => x"49",
   709 => x"c8",
   710 => x"29",
   711 => x"c3",
   712 => x"ff",
   713 => x"99",
   714 => x"73",
   715 => x"09",
   716 => x"97",
   717 => x"79",
   718 => x"09",
   719 => x"d4",
   720 => x"66",
   721 => x"49",
   722 => x"c3",
   723 => x"ff",
   724 => x"99",
   725 => x"73",
   726 => x"09",
   727 => x"97",
   728 => x"79",
   729 => x"09",
   730 => x"d0",
   731 => x"66",
   732 => x"49",
   733 => x"d0",
   734 => x"29",
   735 => x"c3",
   736 => x"ff",
   737 => x"99",
   738 => x"73",
   739 => x"09",
   740 => x"97",
   741 => x"79",
   742 => x"09",
   743 => x"97",
   744 => x"6b",
   745 => x"48",
   746 => x"c4",
   747 => x"a6",
   748 => x"58",
   749 => x"6e",
   750 => x"4c",
   751 => x"c3",
   752 => x"ff",
   753 => x"9c",
   754 => x"c9",
   755 => x"f0",
   756 => x"ff",
   757 => x"4a",
   758 => x"c3",
   759 => x"ff",
   760 => x"ac",
   761 => x"05",
   762 => x"da",
   763 => x"87",
   764 => x"c3",
   765 => x"ff",
   766 => x"97",
   767 => x"7b",
   768 => x"97",
   769 => x"6b",
   770 => x"48",
   771 => x"c4",
   772 => x"a6",
   773 => x"58",
   774 => x"6e",
   775 => x"4c",
   776 => x"c3",
   777 => x"ff",
   778 => x"9c",
   779 => x"c1",
   780 => x"8a",
   781 => x"02",
   782 => x"c6",
   783 => x"87",
   784 => x"c3",
   785 => x"ff",
   786 => x"ac",
   787 => x"02",
   788 => x"e6",
   789 => x"87",
   790 => x"74",
   791 => x"49",
   792 => x"c4",
   793 => x"b7",
   794 => x"29",
   795 => x"c0",
   796 => x"f0",
   797 => x"81",
   798 => x"71",
   799 => x"1e",
   800 => x"c0",
   801 => x"ea",
   802 => x"db",
   803 => x"87",
   804 => x"74",
   805 => x"49",
   806 => x"cf",
   807 => x"99",
   808 => x"c0",
   809 => x"f0",
   810 => x"81",
   811 => x"71",
   812 => x"1e",
   813 => x"c0",
   814 => x"ea",
   815 => x"ce",
   816 => x"87",
   817 => x"74",
   818 => x"48",
   819 => x"f4",
   820 => x"8e",
   821 => x"c2",
   822 => x"87",
   823 => x"26",
   824 => x"4d",
   825 => x"26",
   826 => x"4c",
   827 => x"26",
   828 => x"4b",
   829 => x"26",
   830 => x"4f",
   831 => x"1e",
   832 => x"c0",
   833 => x"49",
   834 => x"c0",
   835 => x"f6",
   836 => x"e4",
   837 => x"c0",
   838 => x"c0",
   839 => x"48",
   840 => x"c3",
   841 => x"ff",
   842 => x"50",
   843 => x"c1",
   844 => x"81",
   845 => x"c3",
   846 => x"c8",
   847 => x"b7",
   848 => x"a9",
   849 => x"04",
   850 => x"ee",
   851 => x"87",
   852 => x"26",
   853 => x"4f",
   854 => x"0e",
   855 => x"5e",
   856 => x"5b",
   857 => x"5c",
   858 => x"0e",
   859 => x"c0",
   860 => x"f6",
   861 => x"e4",
   862 => x"c0",
   863 => x"c0",
   864 => x"4c",
   865 => x"ff",
   866 => x"db",
   867 => x"87",
   868 => x"c4",
   869 => x"f8",
   870 => x"df",
   871 => x"4b",
   872 => x"c0",
   873 => x"1e",
   874 => x"c0",
   875 => x"ff",
   876 => x"f0",
   877 => x"c1",
   878 => x"f7",
   879 => x"1e",
   880 => x"fc",
   881 => x"cf",
   882 => x"87",
   883 => x"c8",
   884 => x"86",
   885 => x"c1",
   886 => x"a8",
   887 => x"05",
   888 => x"c0",
   889 => x"e6",
   890 => x"87",
   891 => x"c3",
   892 => x"ff",
   893 => x"97",
   894 => x"7c",
   895 => x"c1",
   896 => x"c0",
   897 => x"c0",
   898 => x"c0",
   899 => x"c0",
   900 => x"c0",
   901 => x"1e",
   902 => x"c0",
   903 => x"e1",
   904 => x"f0",
   905 => x"c1",
   906 => x"e9",
   907 => x"1e",
   908 => x"fb",
   909 => x"f3",
   910 => x"87",
   911 => x"c8",
   912 => x"86",
   913 => x"70",
   914 => x"98",
   915 => x"05",
   916 => x"c8",
   917 => x"87",
   918 => x"c3",
   919 => x"ff",
   920 => x"97",
   921 => x"7c",
   922 => x"c1",
   923 => x"48",
   924 => x"cb",
   925 => x"87",
   926 => x"fe",
   927 => x"de",
   928 => x"87",
   929 => x"c1",
   930 => x"8b",
   931 => x"05",
   932 => x"ff",
   933 => x"c1",
   934 => x"87",
   935 => x"c0",
   936 => x"48",
   937 => x"fe",
   938 => x"cd",
   939 => x"87",
   940 => x"43",
   941 => x"4d",
   942 => x"44",
   943 => x"34",
   944 => x"31",
   945 => x"20",
   946 => x"25",
   947 => x"64",
   948 => x"0a",
   949 => x"00",
   950 => x"43",
   951 => x"4d",
   952 => x"44",
   953 => x"35",
   954 => x"35",
   955 => x"20",
   956 => x"25",
   957 => x"64",
   958 => x"0a",
   959 => x"00",
   960 => x"43",
   961 => x"4d",
   962 => x"44",
   963 => x"34",
   964 => x"31",
   965 => x"20",
   966 => x"25",
   967 => x"64",
   968 => x"0a",
   969 => x"00",
   970 => x"43",
   971 => x"4d",
   972 => x"44",
   973 => x"35",
   974 => x"35",
   975 => x"20",
   976 => x"25",
   977 => x"64",
   978 => x"0a",
   979 => x"00",
   980 => x"69",
   981 => x"6e",
   982 => x"69",
   983 => x"74",
   984 => x"20",
   985 => x"25",
   986 => x"64",
   987 => x"0a",
   988 => x"20",
   989 => x"20",
   990 => x"00",
   991 => x"69",
   992 => x"6e",
   993 => x"69",
   994 => x"74",
   995 => x"20",
   996 => x"25",
   997 => x"64",
   998 => x"0a",
   999 => x"20",
  1000 => x"20",
  1001 => x"00",
  1002 => x"43",
  1003 => x"6d",
  1004 => x"64",
  1005 => x"5f",
  1006 => x"69",
  1007 => x"6e",
  1008 => x"69",
  1009 => x"74",
  1010 => x"0a",
  1011 => x"00",
  1012 => x"43",
  1013 => x"4d",
  1014 => x"44",
  1015 => x"38",
  1016 => x"5f",
  1017 => x"34",
  1018 => x"20",
  1019 => x"72",
  1020 => x"65",
  1021 => x"73",
  1022 => x"70",
  1023 => x"6f",
  1024 => x"6e",
  1025 => x"73",
  1026 => x"65",
  1027 => x"3a",
  1028 => x"20",
  1029 => x"25",
  1030 => x"64",
  1031 => x"0a",
  1032 => x"00",
  1033 => x"43",
  1034 => x"4d",
  1035 => x"44",
  1036 => x"35",
  1037 => x"38",
  1038 => x"20",
  1039 => x"25",
  1040 => x"64",
  1041 => x"0a",
  1042 => x"20",
  1043 => x"20",
  1044 => x"00",
  1045 => x"43",
  1046 => x"4d",
  1047 => x"44",
  1048 => x"35",
  1049 => x"38",
  1050 => x"5f",
  1051 => x"32",
  1052 => x"20",
  1053 => x"25",
  1054 => x"64",
  1055 => x"0a",
  1056 => x"20",
  1057 => x"20",
  1058 => x"00",
  1059 => x"43",
  1060 => x"4d",
  1061 => x"44",
  1062 => x"35",
  1063 => x"38",
  1064 => x"20",
  1065 => x"25",
  1066 => x"64",
  1067 => x"0a",
  1068 => x"20",
  1069 => x"20",
  1070 => x"00",
  1071 => x"53",
  1072 => x"44",
  1073 => x"48",
  1074 => x"43",
  1075 => x"20",
  1076 => x"49",
  1077 => x"6e",
  1078 => x"69",
  1079 => x"74",
  1080 => x"69",
  1081 => x"61",
  1082 => x"6c",
  1083 => x"69",
  1084 => x"7a",
  1085 => x"61",
  1086 => x"74",
  1087 => x"69",
  1088 => x"6f",
  1089 => x"6e",
  1090 => x"20",
  1091 => x"65",
  1092 => x"72",
  1093 => x"72",
  1094 => x"6f",
  1095 => x"72",
  1096 => x"21",
  1097 => x"0a",
  1098 => x"00",
  1099 => x"63",
  1100 => x"6d",
  1101 => x"64",
  1102 => x"5f",
  1103 => x"43",
  1104 => x"4d",
  1105 => x"44",
  1106 => x"38",
  1107 => x"20",
  1108 => x"72",
  1109 => x"65",
  1110 => x"73",
  1111 => x"70",
  1112 => x"6f",
  1113 => x"6e",
  1114 => x"73",
  1115 => x"65",
  1116 => x"3a",
  1117 => x"20",
  1118 => x"25",
  1119 => x"64",
  1120 => x"0a",
  1121 => x"00",
  1122 => x"52",
  1123 => x"65",
  1124 => x"61",
  1125 => x"64",
  1126 => x"20",
  1127 => x"63",
  1128 => x"6f",
  1129 => x"6d",
  1130 => x"6d",
  1131 => x"61",
  1132 => x"6e",
  1133 => x"64",
  1134 => x"20",
  1135 => x"66",
  1136 => x"61",
  1137 => x"69",
  1138 => x"6c",
  1139 => x"65",
  1140 => x"64",
  1141 => x"20",
  1142 => x"61",
  1143 => x"74",
  1144 => x"20",
  1145 => x"25",
  1146 => x"64",
  1147 => x"20",
  1148 => x"28",
  1149 => x"25",
  1150 => x"64",
  1151 => x"29",
  1152 => x"0a",
  1153 => x"00",
  1154 => x"0e",
  1155 => x"5e",
  1156 => x"5b",
  1157 => x"5c",
  1158 => x"0e",
  1159 => x"c0",
  1160 => x"f6",
  1161 => x"e4",
  1162 => x"c0",
  1163 => x"c0",
  1164 => x"4c",
  1165 => x"c3",
  1166 => x"ff",
  1167 => x"97",
  1168 => x"7c",
  1169 => x"cf",
  1170 => x"ea",
  1171 => x"1e",
  1172 => x"c0",
  1173 => x"e4",
  1174 => x"f4",
  1175 => x"87",
  1176 => x"c4",
  1177 => x"86",
  1178 => x"d3",
  1179 => x"4b",
  1180 => x"c0",
  1181 => x"1e",
  1182 => x"c0",
  1183 => x"ff",
  1184 => x"f0",
  1185 => x"c1",
  1186 => x"c1",
  1187 => x"1e",
  1188 => x"f7",
  1189 => x"db",
  1190 => x"87",
  1191 => x"c8",
  1192 => x"86",
  1193 => x"70",
  1194 => x"98",
  1195 => x"05",
  1196 => x"c8",
  1197 => x"87",
  1198 => x"c3",
  1199 => x"ff",
  1200 => x"97",
  1201 => x"7c",
  1202 => x"c1",
  1203 => x"48",
  1204 => x"cb",
  1205 => x"87",
  1206 => x"fa",
  1207 => x"c6",
  1208 => x"87",
  1209 => x"c1",
  1210 => x"8b",
  1211 => x"05",
  1212 => x"ff",
  1213 => x"dd",
  1214 => x"87",
  1215 => x"c0",
  1216 => x"48",
  1217 => x"f9",
  1218 => x"f5",
  1219 => x"87",
  1220 => x"0e",
  1221 => x"5e",
  1222 => x"5b",
  1223 => x"5c",
  1224 => x"0e",
  1225 => x"1e",
  1226 => x"c0",
  1227 => x"f6",
  1228 => x"e4",
  1229 => x"c0",
  1230 => x"c0",
  1231 => x"4c",
  1232 => x"f9",
  1233 => x"ec",
  1234 => x"87",
  1235 => x"c6",
  1236 => x"ea",
  1237 => x"1e",
  1238 => x"c0",
  1239 => x"e1",
  1240 => x"f0",
  1241 => x"c1",
  1242 => x"c8",
  1243 => x"1e",
  1244 => x"f6",
  1245 => x"e3",
  1246 => x"87",
  1247 => x"70",
  1248 => x"4b",
  1249 => x"73",
  1250 => x"1e",
  1251 => x"d1",
  1252 => x"cb",
  1253 => x"1e",
  1254 => x"c0",
  1255 => x"f2",
  1256 => x"e3",
  1257 => x"87",
  1258 => x"d0",
  1259 => x"86",
  1260 => x"c1",
  1261 => x"ab",
  1262 => x"02",
  1263 => x"c8",
  1264 => x"87",
  1265 => x"fe",
  1266 => x"ce",
  1267 => x"87",
  1268 => x"c0",
  1269 => x"48",
  1270 => x"c1",
  1271 => x"f0",
  1272 => x"87",
  1273 => x"f4",
  1274 => x"e3",
  1275 => x"87",
  1276 => x"70",
  1277 => x"49",
  1278 => x"cf",
  1279 => x"ff",
  1280 => x"ff",
  1281 => x"99",
  1282 => x"c6",
  1283 => x"ea",
  1284 => x"a9",
  1285 => x"02",
  1286 => x"c8",
  1287 => x"87",
  1288 => x"fd",
  1289 => x"f7",
  1290 => x"87",
  1291 => x"c0",
  1292 => x"48",
  1293 => x"c1",
  1294 => x"d9",
  1295 => x"87",
  1296 => x"c3",
  1297 => x"ff",
  1298 => x"97",
  1299 => x"7c",
  1300 => x"c0",
  1301 => x"f1",
  1302 => x"4b",
  1303 => x"f8",
  1304 => x"fc",
  1305 => x"87",
  1306 => x"70",
  1307 => x"98",
  1308 => x"02",
  1309 => x"c0",
  1310 => x"f8",
  1311 => x"87",
  1312 => x"c0",
  1313 => x"1e",
  1314 => x"c0",
  1315 => x"ff",
  1316 => x"f0",
  1317 => x"c1",
  1318 => x"fa",
  1319 => x"1e",
  1320 => x"f5",
  1321 => x"d7",
  1322 => x"87",
  1323 => x"c8",
  1324 => x"86",
  1325 => x"70",
  1326 => x"98",
  1327 => x"05",
  1328 => x"c0",
  1329 => x"e5",
  1330 => x"87",
  1331 => x"c3",
  1332 => x"ff",
  1333 => x"97",
  1334 => x"7c",
  1335 => x"97",
  1336 => x"6c",
  1337 => x"48",
  1338 => x"c4",
  1339 => x"a6",
  1340 => x"58",
  1341 => x"6e",
  1342 => x"49",
  1343 => x"c3",
  1344 => x"ff",
  1345 => x"99",
  1346 => x"97",
  1347 => x"7c",
  1348 => x"97",
  1349 => x"7c",
  1350 => x"97",
  1351 => x"7c",
  1352 => x"97",
  1353 => x"7c",
  1354 => x"c1",
  1355 => x"c0",
  1356 => x"99",
  1357 => x"02",
  1358 => x"c4",
  1359 => x"87",
  1360 => x"c1",
  1361 => x"48",
  1362 => x"d5",
  1363 => x"87",
  1364 => x"c0",
  1365 => x"48",
  1366 => x"d1",
  1367 => x"87",
  1368 => x"c2",
  1369 => x"ab",
  1370 => x"05",
  1371 => x"c4",
  1372 => x"87",
  1373 => x"c0",
  1374 => x"48",
  1375 => x"c8",
  1376 => x"87",
  1377 => x"c1",
  1378 => x"8b",
  1379 => x"05",
  1380 => x"fe",
  1381 => x"f0",
  1382 => x"87",
  1383 => x"c0",
  1384 => x"48",
  1385 => x"26",
  1386 => x"f7",
  1387 => x"cc",
  1388 => x"87",
  1389 => x"0e",
  1390 => x"5e",
  1391 => x"5b",
  1392 => x"5c",
  1393 => x"5d",
  1394 => x"0e",
  1395 => x"c0",
  1396 => x"f6",
  1397 => x"e4",
  1398 => x"c0",
  1399 => x"c0",
  1400 => x"4c",
  1401 => x"48",
  1402 => x"c4",
  1403 => x"a0",
  1404 => x"4b",
  1405 => x"c1",
  1406 => x"c8",
  1407 => x"e8",
  1408 => x"48",
  1409 => x"c1",
  1410 => x"78",
  1411 => x"c0",
  1412 => x"f6",
  1413 => x"e4",
  1414 => x"c0",
  1415 => x"c8",
  1416 => x"48",
  1417 => x"c0",
  1418 => x"e0",
  1419 => x"50",
  1420 => x"c7",
  1421 => x"4d",
  1422 => x"c3",
  1423 => x"97",
  1424 => x"7b",
  1425 => x"f6",
  1426 => x"eb",
  1427 => x"87",
  1428 => x"c2",
  1429 => x"97",
  1430 => x"7b",
  1431 => x"c3",
  1432 => x"ff",
  1433 => x"97",
  1434 => x"7c",
  1435 => x"c0",
  1436 => x"1e",
  1437 => x"c0",
  1438 => x"e5",
  1439 => x"d0",
  1440 => x"c1",
  1441 => x"c0",
  1442 => x"1e",
  1443 => x"f3",
  1444 => x"dc",
  1445 => x"87",
  1446 => x"c8",
  1447 => x"86",
  1448 => x"c1",
  1449 => x"a8",
  1450 => x"05",
  1451 => x"c2",
  1452 => x"87",
  1453 => x"c1",
  1454 => x"4d",
  1455 => x"c2",
  1456 => x"ad",
  1457 => x"05",
  1458 => x"c5",
  1459 => x"87",
  1460 => x"c0",
  1461 => x"48",
  1462 => x"c0",
  1463 => x"ec",
  1464 => x"87",
  1465 => x"c1",
  1466 => x"8d",
  1467 => x"05",
  1468 => x"ff",
  1469 => x"cf",
  1470 => x"87",
  1471 => x"fc",
  1472 => x"c2",
  1473 => x"87",
  1474 => x"c1",
  1475 => x"c8",
  1476 => x"ec",
  1477 => x"58",
  1478 => x"c1",
  1479 => x"c8",
  1480 => x"e8",
  1481 => x"bf",
  1482 => x"05",
  1483 => x"cd",
  1484 => x"87",
  1485 => x"c1",
  1486 => x"1e",
  1487 => x"c0",
  1488 => x"ff",
  1489 => x"f0",
  1490 => x"c1",
  1491 => x"d0",
  1492 => x"1e",
  1493 => x"f2",
  1494 => x"ea",
  1495 => x"87",
  1496 => x"c8",
  1497 => x"86",
  1498 => x"c3",
  1499 => x"ff",
  1500 => x"97",
  1501 => x"7c",
  1502 => x"c3",
  1503 => x"53",
  1504 => x"c3",
  1505 => x"ff",
  1506 => x"54",
  1507 => x"c1",
  1508 => x"48",
  1509 => x"f5",
  1510 => x"cf",
  1511 => x"87",
  1512 => x"0e",
  1513 => x"5e",
  1514 => x"5b",
  1515 => x"5c",
  1516 => x"5d",
  1517 => x"0e",
  1518 => x"1e",
  1519 => x"c0",
  1520 => x"f6",
  1521 => x"e4",
  1522 => x"c0",
  1523 => x"c0",
  1524 => x"4b",
  1525 => x"c0",
  1526 => x"4d",
  1527 => x"c3",
  1528 => x"ff",
  1529 => x"97",
  1530 => x"7b",
  1531 => x"c0",
  1532 => x"f6",
  1533 => x"e4",
  1534 => x"c0",
  1535 => x"c4",
  1536 => x"48",
  1537 => x"c2",
  1538 => x"50",
  1539 => x"c0",
  1540 => x"f6",
  1541 => x"e4",
  1542 => x"c0",
  1543 => x"c8",
  1544 => x"48",
  1545 => x"c1",
  1546 => x"50",
  1547 => x"c3",
  1548 => x"ff",
  1549 => x"97",
  1550 => x"7b",
  1551 => x"d4",
  1552 => x"66",
  1553 => x"1e",
  1554 => x"c0",
  1555 => x"ff",
  1556 => x"f0",
  1557 => x"c1",
  1558 => x"d1",
  1559 => x"1e",
  1560 => x"f1",
  1561 => x"e7",
  1562 => x"87",
  1563 => x"c8",
  1564 => x"86",
  1565 => x"70",
  1566 => x"98",
  1567 => x"05",
  1568 => x"c1",
  1569 => x"c9",
  1570 => x"87",
  1571 => x"c5",
  1572 => x"ee",
  1573 => x"cd",
  1574 => x"df",
  1575 => x"4a",
  1576 => x"c3",
  1577 => x"ff",
  1578 => x"97",
  1579 => x"7b",
  1580 => x"97",
  1581 => x"6b",
  1582 => x"48",
  1583 => x"c4",
  1584 => x"a6",
  1585 => x"58",
  1586 => x"6e",
  1587 => x"49",
  1588 => x"c3",
  1589 => x"ff",
  1590 => x"99",
  1591 => x"c3",
  1592 => x"fe",
  1593 => x"a9",
  1594 => x"05",
  1595 => x"de",
  1596 => x"87",
  1597 => x"c0",
  1598 => x"4c",
  1599 => x"ef",
  1600 => x"dd",
  1601 => x"87",
  1602 => x"d8",
  1603 => x"66",
  1604 => x"08",
  1605 => x"78",
  1606 => x"08",
  1607 => x"d8",
  1608 => x"66",
  1609 => x"48",
  1610 => x"c4",
  1611 => x"80",
  1612 => x"dc",
  1613 => x"a6",
  1614 => x"58",
  1615 => x"c1",
  1616 => x"84",
  1617 => x"c2",
  1618 => x"c0",
  1619 => x"b7",
  1620 => x"ac",
  1621 => x"04",
  1622 => x"e7",
  1623 => x"87",
  1624 => x"c1",
  1625 => x"4a",
  1626 => x"4d",
  1627 => x"c1",
  1628 => x"8a",
  1629 => x"05",
  1630 => x"ff",
  1631 => x"c7",
  1632 => x"87",
  1633 => x"c3",
  1634 => x"ff",
  1635 => x"53",
  1636 => x"c0",
  1637 => x"f6",
  1638 => x"e4",
  1639 => x"c0",
  1640 => x"c4",
  1641 => x"48",
  1642 => x"c3",
  1643 => x"50",
  1644 => x"75",
  1645 => x"48",
  1646 => x"26",
  1647 => x"f3",
  1648 => x"c5",
  1649 => x"87",
  1650 => x"1e",
  1651 => x"c4",
  1652 => x"66",
  1653 => x"49",
  1654 => x"d8",
  1655 => x"29",
  1656 => x"c3",
  1657 => x"ff",
  1658 => x"99",
  1659 => x"c4",
  1660 => x"66",
  1661 => x"4a",
  1662 => x"c8",
  1663 => x"2a",
  1664 => x"cf",
  1665 => x"fc",
  1666 => x"c0",
  1667 => x"9a",
  1668 => x"72",
  1669 => x"b1",
  1670 => x"c4",
  1671 => x"66",
  1672 => x"4a",
  1673 => x"c8",
  1674 => x"32",
  1675 => x"c0",
  1676 => x"ff",
  1677 => x"f0",
  1678 => x"c0",
  1679 => x"c0",
  1680 => x"9a",
  1681 => x"72",
  1682 => x"b1",
  1683 => x"c4",
  1684 => x"66",
  1685 => x"4a",
  1686 => x"d8",
  1687 => x"32",
  1688 => x"ff",
  1689 => x"c0",
  1690 => x"c0",
  1691 => x"c0",
  1692 => x"c0",
  1693 => x"9a",
  1694 => x"72",
  1695 => x"b1",
  1696 => x"71",
  1697 => x"48",
  1698 => x"26",
  1699 => x"4f",
  1700 => x"1e",
  1701 => x"c4",
  1702 => x"66",
  1703 => x"49",
  1704 => x"c8",
  1705 => x"29",
  1706 => x"c3",
  1707 => x"ff",
  1708 => x"99",
  1709 => x"c4",
  1710 => x"66",
  1711 => x"4a",
  1712 => x"c8",
  1713 => x"32",
  1714 => x"cf",
  1715 => x"fc",
  1716 => x"c0",
  1717 => x"9a",
  1718 => x"72",
  1719 => x"b1",
  1720 => x"71",
  1721 => x"48",
  1722 => x"26",
  1723 => x"4f",
  1724 => x"1e",
  1725 => x"73",
  1726 => x"1e",
  1727 => x"c0",
  1728 => x"4b",
  1729 => x"d0",
  1730 => x"66",
  1731 => x"48",
  1732 => x"c0",
  1733 => x"b7",
  1734 => x"a8",
  1735 => x"06",
  1736 => x"c0",
  1737 => x"ee",
  1738 => x"87",
  1739 => x"c8",
  1740 => x"66",
  1741 => x"97",
  1742 => x"bf",
  1743 => x"4a",
  1744 => x"c8",
  1745 => x"66",
  1746 => x"48",
  1747 => x"c1",
  1748 => x"80",
  1749 => x"cc",
  1750 => x"a6",
  1751 => x"58",
  1752 => x"cc",
  1753 => x"66",
  1754 => x"97",
  1755 => x"bf",
  1756 => x"49",
  1757 => x"cc",
  1758 => x"66",
  1759 => x"48",
  1760 => x"c1",
  1761 => x"80",
  1762 => x"d0",
  1763 => x"a6",
  1764 => x"58",
  1765 => x"71",
  1766 => x"b7",
  1767 => x"aa",
  1768 => x"02",
  1769 => x"c4",
  1770 => x"87",
  1771 => x"c1",
  1772 => x"48",
  1773 => x"cc",
  1774 => x"87",
  1775 => x"c1",
  1776 => x"83",
  1777 => x"d0",
  1778 => x"66",
  1779 => x"b7",
  1780 => x"ab",
  1781 => x"04",
  1782 => x"ff",
  1783 => x"d2",
  1784 => x"87",
  1785 => x"c0",
  1786 => x"48",
  1787 => x"c4",
  1788 => x"87",
  1789 => x"26",
  1790 => x"4d",
  1791 => x"26",
  1792 => x"4c",
  1793 => x"26",
  1794 => x"4b",
  1795 => x"26",
  1796 => x"4f",
  1797 => x"0e",
  1798 => x"5e",
  1799 => x"5b",
  1800 => x"5c",
  1801 => x"5d",
  1802 => x"0e",
  1803 => x"c1",
  1804 => x"d1",
  1805 => x"ea",
  1806 => x"48",
  1807 => x"ff",
  1808 => x"78",
  1809 => x"c1",
  1810 => x"d0",
  1811 => x"fa",
  1812 => x"48",
  1813 => x"c0",
  1814 => x"78",
  1815 => x"c0",
  1816 => x"ea",
  1817 => x"c0",
  1818 => x"1e",
  1819 => x"da",
  1820 => x"ee",
  1821 => x"87",
  1822 => x"c1",
  1823 => x"c8",
  1824 => x"f2",
  1825 => x"1e",
  1826 => x"c0",
  1827 => x"1e",
  1828 => x"fb",
  1829 => x"c1",
  1830 => x"87",
  1831 => x"cc",
  1832 => x"86",
  1833 => x"70",
  1834 => x"98",
  1835 => x"05",
  1836 => x"c5",
  1837 => x"87",
  1838 => x"c0",
  1839 => x"48",
  1840 => x"cb",
  1841 => x"c7",
  1842 => x"87",
  1843 => x"c0",
  1844 => x"4b",
  1845 => x"c1",
  1846 => x"d1",
  1847 => x"e6",
  1848 => x"48",
  1849 => x"c1",
  1850 => x"78",
  1851 => x"c8",
  1852 => x"1e",
  1853 => x"c0",
  1854 => x"ea",
  1855 => x"cd",
  1856 => x"1e",
  1857 => x"c1",
  1858 => x"c9",
  1859 => x"e8",
  1860 => x"1e",
  1861 => x"fd",
  1862 => x"f4",
  1863 => x"87",
  1864 => x"cc",
  1865 => x"86",
  1866 => x"70",
  1867 => x"98",
  1868 => x"05",
  1869 => x"c6",
  1870 => x"87",
  1871 => x"c1",
  1872 => x"d1",
  1873 => x"e6",
  1874 => x"48",
  1875 => x"c0",
  1876 => x"78",
  1877 => x"c8",
  1878 => x"1e",
  1879 => x"c0",
  1880 => x"ea",
  1881 => x"d6",
  1882 => x"1e",
  1883 => x"c1",
  1884 => x"ca",
  1885 => x"c4",
  1886 => x"1e",
  1887 => x"fd",
  1888 => x"da",
  1889 => x"87",
  1890 => x"cc",
  1891 => x"86",
  1892 => x"70",
  1893 => x"98",
  1894 => x"05",
  1895 => x"c6",
  1896 => x"87",
  1897 => x"c1",
  1898 => x"d1",
  1899 => x"e6",
  1900 => x"48",
  1901 => x"c0",
  1902 => x"78",
  1903 => x"c8",
  1904 => x"1e",
  1905 => x"c0",
  1906 => x"ea",
  1907 => x"df",
  1908 => x"1e",
  1909 => x"c1",
  1910 => x"ca",
  1911 => x"c4",
  1912 => x"1e",
  1913 => x"fd",
  1914 => x"c0",
  1915 => x"87",
  1916 => x"cc",
  1917 => x"86",
  1918 => x"70",
  1919 => x"98",
  1920 => x"05",
  1921 => x"c5",
  1922 => x"87",
  1923 => x"c0",
  1924 => x"48",
  1925 => x"c9",
  1926 => x"f2",
  1927 => x"87",
  1928 => x"c1",
  1929 => x"d1",
  1930 => x"e6",
  1931 => x"bf",
  1932 => x"1e",
  1933 => x"c0",
  1934 => x"ea",
  1935 => x"e8",
  1936 => x"1e",
  1937 => x"c0",
  1938 => x"e7",
  1939 => x"f8",
  1940 => x"87",
  1941 => x"c8",
  1942 => x"86",
  1943 => x"c1",
  1944 => x"d1",
  1945 => x"e6",
  1946 => x"bf",
  1947 => x"02",
  1948 => x"c1",
  1949 => x"fa",
  1950 => x"87",
  1951 => x"c1",
  1952 => x"c8",
  1953 => x"f2",
  1954 => x"4d",
  1955 => x"48",
  1956 => x"c6",
  1957 => x"fe",
  1958 => x"a0",
  1959 => x"4c",
  1960 => x"c8",
  1961 => x"c0",
  1962 => x"1e",
  1963 => x"70",
  1964 => x"1e",
  1965 => x"da",
  1966 => x"f3",
  1967 => x"87",
  1968 => x"c8",
  1969 => x"86",
  1970 => x"c8",
  1971 => x"a4",
  1972 => x"49",
  1973 => x"69",
  1974 => x"4b",
  1975 => x"c1",
  1976 => x"d0",
  1977 => x"f0",
  1978 => x"9f",
  1979 => x"bf",
  1980 => x"49",
  1981 => x"c5",
  1982 => x"d6",
  1983 => x"ea",
  1984 => x"a9",
  1985 => x"05",
  1986 => x"c0",
  1987 => x"ce",
  1988 => x"87",
  1989 => x"c8",
  1990 => x"a4",
  1991 => x"49",
  1992 => x"69",
  1993 => x"1e",
  1994 => x"fa",
  1995 => x"e5",
  1996 => x"87",
  1997 => x"c4",
  1998 => x"86",
  1999 => x"70",
  2000 => x"4b",
  2001 => x"dd",
  2002 => x"87",
  2003 => x"c7",
  2004 => x"fe",
  2005 => x"a5",
  2006 => x"49",
  2007 => x"9f",
  2008 => x"69",
  2009 => x"49",
  2010 => x"ca",
  2011 => x"e9",
  2012 => x"d5",
  2013 => x"a9",
  2014 => x"02",
  2015 => x"c0",
  2016 => x"ce",
  2017 => x"87",
  2018 => x"c0",
  2019 => x"e7",
  2020 => x"fd",
  2021 => x"1e",
  2022 => x"d7",
  2023 => x"e3",
  2024 => x"87",
  2025 => x"c4",
  2026 => x"86",
  2027 => x"c0",
  2028 => x"48",
  2029 => x"c8",
  2030 => x"ca",
  2031 => x"87",
  2032 => x"73",
  2033 => x"1e",
  2034 => x"c0",
  2035 => x"e8",
  2036 => x"db",
  2037 => x"1e",
  2038 => x"c0",
  2039 => x"e6",
  2040 => x"d3",
  2041 => x"87",
  2042 => x"c1",
  2043 => x"c8",
  2044 => x"f2",
  2045 => x"1e",
  2046 => x"73",
  2047 => x"1e",
  2048 => x"f7",
  2049 => x"e5",
  2050 => x"87",
  2051 => x"d0",
  2052 => x"86",
  2053 => x"70",
  2054 => x"98",
  2055 => x"05",
  2056 => x"c0",
  2057 => x"c5",
  2058 => x"87",
  2059 => x"c0",
  2060 => x"48",
  2061 => x"c7",
  2062 => x"ea",
  2063 => x"87",
  2064 => x"c0",
  2065 => x"e8",
  2066 => x"f3",
  2067 => x"1e",
  2068 => x"d6",
  2069 => x"f5",
  2070 => x"87",
  2071 => x"c4",
  2072 => x"86",
  2073 => x"c8",
  2074 => x"c0",
  2075 => x"1e",
  2076 => x"c1",
  2077 => x"c8",
  2078 => x"f2",
  2079 => x"1e",
  2080 => x"d9",
  2081 => x"c0",
  2082 => x"87",
  2083 => x"c0",
  2084 => x"ea",
  2085 => x"fb",
  2086 => x"1e",
  2087 => x"c0",
  2088 => x"e5",
  2089 => x"e2",
  2090 => x"87",
  2091 => x"c8",
  2092 => x"1e",
  2093 => x"c0",
  2094 => x"eb",
  2095 => x"d3",
  2096 => x"1e",
  2097 => x"c1",
  2098 => x"ca",
  2099 => x"c4",
  2100 => x"1e",
  2101 => x"fa",
  2102 => x"c4",
  2103 => x"87",
  2104 => x"d8",
  2105 => x"86",
  2106 => x"70",
  2107 => x"98",
  2108 => x"05",
  2109 => x"c0",
  2110 => x"c9",
  2111 => x"87",
  2112 => x"c1",
  2113 => x"d0",
  2114 => x"fa",
  2115 => x"48",
  2116 => x"c1",
  2117 => x"78",
  2118 => x"c0",
  2119 => x"e4",
  2120 => x"87",
  2121 => x"c8",
  2122 => x"1e",
  2123 => x"c0",
  2124 => x"eb",
  2125 => x"dc",
  2126 => x"1e",
  2127 => x"c1",
  2128 => x"c9",
  2129 => x"e8",
  2130 => x"1e",
  2131 => x"f9",
  2132 => x"e6",
  2133 => x"87",
  2134 => x"cc",
  2135 => x"86",
  2136 => x"70",
  2137 => x"98",
  2138 => x"02",
  2139 => x"c0",
  2140 => x"cf",
  2141 => x"87",
  2142 => x"c0",
  2143 => x"e9",
  2144 => x"da",
  2145 => x"1e",
  2146 => x"c0",
  2147 => x"e4",
  2148 => x"e7",
  2149 => x"87",
  2150 => x"c4",
  2151 => x"86",
  2152 => x"c0",
  2153 => x"48",
  2154 => x"c6",
  2155 => x"cd",
  2156 => x"87",
  2157 => x"c1",
  2158 => x"d0",
  2159 => x"f0",
  2160 => x"97",
  2161 => x"bf",
  2162 => x"49",
  2163 => x"c1",
  2164 => x"d5",
  2165 => x"a9",
  2166 => x"05",
  2167 => x"c0",
  2168 => x"cd",
  2169 => x"87",
  2170 => x"c1",
  2171 => x"d0",
  2172 => x"f1",
  2173 => x"97",
  2174 => x"bf",
  2175 => x"49",
  2176 => x"c2",
  2177 => x"ea",
  2178 => x"a9",
  2179 => x"02",
  2180 => x"c0",
  2181 => x"c5",
  2182 => x"87",
  2183 => x"c0",
  2184 => x"48",
  2185 => x"c5",
  2186 => x"ee",
  2187 => x"87",
  2188 => x"c1",
  2189 => x"c8",
  2190 => x"f2",
  2191 => x"97",
  2192 => x"bf",
  2193 => x"49",
  2194 => x"c3",
  2195 => x"e9",
  2196 => x"a9",
  2197 => x"02",
  2198 => x"c0",
  2199 => x"d2",
  2200 => x"87",
  2201 => x"c1",
  2202 => x"c8",
  2203 => x"f2",
  2204 => x"97",
  2205 => x"bf",
  2206 => x"49",
  2207 => x"c3",
  2208 => x"eb",
  2209 => x"a9",
  2210 => x"02",
  2211 => x"c0",
  2212 => x"c5",
  2213 => x"87",
  2214 => x"c0",
  2215 => x"48",
  2216 => x"c5",
  2217 => x"cf",
  2218 => x"87",
  2219 => x"c1",
  2220 => x"c8",
  2221 => x"fd",
  2222 => x"97",
  2223 => x"bf",
  2224 => x"49",
  2225 => x"71",
  2226 => x"99",
  2227 => x"05",
  2228 => x"c0",
  2229 => x"cc",
  2230 => x"87",
  2231 => x"c1",
  2232 => x"c8",
  2233 => x"fe",
  2234 => x"97",
  2235 => x"bf",
  2236 => x"49",
  2237 => x"c2",
  2238 => x"a9",
  2239 => x"02",
  2240 => x"c0",
  2241 => x"c5",
  2242 => x"87",
  2243 => x"c0",
  2244 => x"48",
  2245 => x"c4",
  2246 => x"f2",
  2247 => x"87",
  2248 => x"c1",
  2249 => x"c8",
  2250 => x"ff",
  2251 => x"97",
  2252 => x"bf",
  2253 => x"48",
  2254 => x"c1",
  2255 => x"d0",
  2256 => x"f6",
  2257 => x"58",
  2258 => x"c1",
  2259 => x"d0",
  2260 => x"f2",
  2261 => x"bf",
  2262 => x"48",
  2263 => x"c1",
  2264 => x"88",
  2265 => x"c1",
  2266 => x"d0",
  2267 => x"fa",
  2268 => x"58",
  2269 => x"c1",
  2270 => x"c9",
  2271 => x"c0",
  2272 => x"97",
  2273 => x"bf",
  2274 => x"49",
  2275 => x"73",
  2276 => x"81",
  2277 => x"c1",
  2278 => x"c9",
  2279 => x"c1",
  2280 => x"97",
  2281 => x"bf",
  2282 => x"4a",
  2283 => x"c8",
  2284 => x"32",
  2285 => x"c1",
  2286 => x"d1",
  2287 => x"c6",
  2288 => x"48",
  2289 => x"72",
  2290 => x"a1",
  2291 => x"78",
  2292 => x"c1",
  2293 => x"c9",
  2294 => x"c2",
  2295 => x"97",
  2296 => x"bf",
  2297 => x"48",
  2298 => x"c1",
  2299 => x"d1",
  2300 => x"de",
  2301 => x"58",
  2302 => x"c1",
  2303 => x"d0",
  2304 => x"fa",
  2305 => x"bf",
  2306 => x"02",
  2307 => x"c2",
  2308 => x"e2",
  2309 => x"87",
  2310 => x"c8",
  2311 => x"1e",
  2312 => x"c0",
  2313 => x"e9",
  2314 => x"f7",
  2315 => x"1e",
  2316 => x"c1",
  2317 => x"ca",
  2318 => x"c4",
  2319 => x"1e",
  2320 => x"f6",
  2321 => x"e9",
  2322 => x"87",
  2323 => x"cc",
  2324 => x"86",
  2325 => x"70",
  2326 => x"98",
  2327 => x"02",
  2328 => x"c0",
  2329 => x"c5",
  2330 => x"87",
  2331 => x"c0",
  2332 => x"48",
  2333 => x"c3",
  2334 => x"da",
  2335 => x"87",
  2336 => x"c1",
  2337 => x"d0",
  2338 => x"f2",
  2339 => x"bf",
  2340 => x"48",
  2341 => x"c4",
  2342 => x"30",
  2343 => x"c1",
  2344 => x"d1",
  2345 => x"e2",
  2346 => x"58",
  2347 => x"c1",
  2348 => x"d0",
  2349 => x"f2",
  2350 => x"bf",
  2351 => x"4a",
  2352 => x"c1",
  2353 => x"d1",
  2354 => x"da",
  2355 => x"5a",
  2356 => x"c1",
  2357 => x"c9",
  2358 => x"d7",
  2359 => x"97",
  2360 => x"bf",
  2361 => x"49",
  2362 => x"c8",
  2363 => x"31",
  2364 => x"c1",
  2365 => x"c9",
  2366 => x"d6",
  2367 => x"97",
  2368 => x"bf",
  2369 => x"4b",
  2370 => x"73",
  2371 => x"a1",
  2372 => x"49",
  2373 => x"c1",
  2374 => x"c9",
  2375 => x"d8",
  2376 => x"97",
  2377 => x"bf",
  2378 => x"4b",
  2379 => x"d0",
  2380 => x"33",
  2381 => x"73",
  2382 => x"a1",
  2383 => x"49",
  2384 => x"c1",
  2385 => x"c9",
  2386 => x"d9",
  2387 => x"97",
  2388 => x"bf",
  2389 => x"4b",
  2390 => x"d8",
  2391 => x"33",
  2392 => x"73",
  2393 => x"a1",
  2394 => x"49",
  2395 => x"c1",
  2396 => x"d1",
  2397 => x"e6",
  2398 => x"59",
  2399 => x"c1",
  2400 => x"d1",
  2401 => x"da",
  2402 => x"bf",
  2403 => x"91",
  2404 => x"c1",
  2405 => x"d1",
  2406 => x"c6",
  2407 => x"bf",
  2408 => x"81",
  2409 => x"c1",
  2410 => x"d1",
  2411 => x"ce",
  2412 => x"59",
  2413 => x"c1",
  2414 => x"c9",
  2415 => x"df",
  2416 => x"97",
  2417 => x"bf",
  2418 => x"4b",
  2419 => x"c8",
  2420 => x"33",
  2421 => x"c1",
  2422 => x"c9",
  2423 => x"de",
  2424 => x"97",
  2425 => x"bf",
  2426 => x"4c",
  2427 => x"74",
  2428 => x"a3",
  2429 => x"4b",
  2430 => x"c1",
  2431 => x"c9",
  2432 => x"e0",
  2433 => x"97",
  2434 => x"bf",
  2435 => x"4c",
  2436 => x"d0",
  2437 => x"34",
  2438 => x"74",
  2439 => x"a3",
  2440 => x"4b",
  2441 => x"c1",
  2442 => x"c9",
  2443 => x"e1",
  2444 => x"97",
  2445 => x"bf",
  2446 => x"4c",
  2447 => x"cf",
  2448 => x"9c",
  2449 => x"d8",
  2450 => x"34",
  2451 => x"74",
  2452 => x"a3",
  2453 => x"4b",
  2454 => x"c1",
  2455 => x"d1",
  2456 => x"d2",
  2457 => x"5b",
  2458 => x"c2",
  2459 => x"8b",
  2460 => x"73",
  2461 => x"92",
  2462 => x"c1",
  2463 => x"d1",
  2464 => x"d2",
  2465 => x"48",
  2466 => x"72",
  2467 => x"a1",
  2468 => x"78",
  2469 => x"c1",
  2470 => x"d0",
  2471 => x"87",
  2472 => x"c1",
  2473 => x"c9",
  2474 => x"c4",
  2475 => x"97",
  2476 => x"bf",
  2477 => x"49",
  2478 => x"c8",
  2479 => x"31",
  2480 => x"c1",
  2481 => x"c9",
  2482 => x"c3",
  2483 => x"97",
  2484 => x"bf",
  2485 => x"4a",
  2486 => x"72",
  2487 => x"a1",
  2488 => x"49",
  2489 => x"c1",
  2490 => x"d1",
  2491 => x"e2",
  2492 => x"59",
  2493 => x"c5",
  2494 => x"31",
  2495 => x"c7",
  2496 => x"ff",
  2497 => x"81",
  2498 => x"c9",
  2499 => x"29",
  2500 => x"c1",
  2501 => x"d1",
  2502 => x"da",
  2503 => x"59",
  2504 => x"c1",
  2505 => x"c9",
  2506 => x"c9",
  2507 => x"97",
  2508 => x"bf",
  2509 => x"4a",
  2510 => x"c8",
  2511 => x"32",
  2512 => x"c1",
  2513 => x"c9",
  2514 => x"c8",
  2515 => x"97",
  2516 => x"bf",
  2517 => x"4b",
  2518 => x"73",
  2519 => x"a2",
  2520 => x"4a",
  2521 => x"c1",
  2522 => x"d1",
  2523 => x"e6",
  2524 => x"5a",
  2525 => x"c1",
  2526 => x"d1",
  2527 => x"da",
  2528 => x"bf",
  2529 => x"92",
  2530 => x"c1",
  2531 => x"d1",
  2532 => x"c6",
  2533 => x"bf",
  2534 => x"82",
  2535 => x"c1",
  2536 => x"d1",
  2537 => x"d6",
  2538 => x"5a",
  2539 => x"c1",
  2540 => x"d1",
  2541 => x"ce",
  2542 => x"48",
  2543 => x"c0",
  2544 => x"78",
  2545 => x"c1",
  2546 => x"d1",
  2547 => x"ca",
  2548 => x"48",
  2549 => x"72",
  2550 => x"a1",
  2551 => x"78",
  2552 => x"c1",
  2553 => x"48",
  2554 => x"f4",
  2555 => x"c0",
  2556 => x"87",
  2557 => x"4e",
  2558 => x"6f",
  2559 => x"20",
  2560 => x"70",
  2561 => x"61",
  2562 => x"72",
  2563 => x"74",
  2564 => x"69",
  2565 => x"74",
  2566 => x"69",
  2567 => x"6f",
  2568 => x"6e",
  2569 => x"20",
  2570 => x"73",
  2571 => x"69",
  2572 => x"67",
  2573 => x"6e",
  2574 => x"61",
  2575 => x"74",
  2576 => x"75",
  2577 => x"72",
  2578 => x"65",
  2579 => x"20",
  2580 => x"66",
  2581 => x"6f",
  2582 => x"75",
  2583 => x"6e",
  2584 => x"64",
  2585 => x"0a",
  2586 => x"00",
  2587 => x"52",
  2588 => x"65",
  2589 => x"61",
  2590 => x"64",
  2591 => x"69",
  2592 => x"6e",
  2593 => x"67",
  2594 => x"20",
  2595 => x"62",
  2596 => x"6f",
  2597 => x"6f",
  2598 => x"74",
  2599 => x"20",
  2600 => x"73",
  2601 => x"65",
  2602 => x"63",
  2603 => x"74",
  2604 => x"6f",
  2605 => x"72",
  2606 => x"20",
  2607 => x"25",
  2608 => x"64",
  2609 => x"0a",
  2610 => x"00",
  2611 => x"52",
  2612 => x"65",
  2613 => x"61",
  2614 => x"64",
  2615 => x"20",
  2616 => x"62",
  2617 => x"6f",
  2618 => x"6f",
  2619 => x"74",
  2620 => x"20",
  2621 => x"73",
  2622 => x"65",
  2623 => x"63",
  2624 => x"74",
  2625 => x"6f",
  2626 => x"72",
  2627 => x"20",
  2628 => x"66",
  2629 => x"72",
  2630 => x"6f",
  2631 => x"6d",
  2632 => x"20",
  2633 => x"66",
  2634 => x"69",
  2635 => x"72",
  2636 => x"73",
  2637 => x"74",
  2638 => x"20",
  2639 => x"70",
  2640 => x"61",
  2641 => x"72",
  2642 => x"74",
  2643 => x"69",
  2644 => x"74",
  2645 => x"69",
  2646 => x"6f",
  2647 => x"6e",
  2648 => x"0a",
  2649 => x"00",
  2650 => x"55",
  2651 => x"6e",
  2652 => x"73",
  2653 => x"75",
  2654 => x"70",
  2655 => x"70",
  2656 => x"6f",
  2657 => x"72",
  2658 => x"74",
  2659 => x"65",
  2660 => x"64",
  2661 => x"20",
  2662 => x"70",
  2663 => x"61",
  2664 => x"72",
  2665 => x"74",
  2666 => x"69",
  2667 => x"74",
  2668 => x"69",
  2669 => x"6f",
  2670 => x"6e",
  2671 => x"20",
  2672 => x"74",
  2673 => x"79",
  2674 => x"70",
  2675 => x"65",
  2676 => x"21",
  2677 => x"0d",
  2678 => x"00",
  2679 => x"46",
  2680 => x"41",
  2681 => x"54",
  2682 => x"33",
  2683 => x"32",
  2684 => x"20",
  2685 => x"20",
  2686 => x"20",
  2687 => x"00",
  2688 => x"52",
  2689 => x"65",
  2690 => x"61",
  2691 => x"64",
  2692 => x"69",
  2693 => x"6e",
  2694 => x"67",
  2695 => x"20",
  2696 => x"4d",
  2697 => x"42",
  2698 => x"52",
  2699 => x"0a",
  2700 => x"00",
  2701 => x"46",
  2702 => x"41",
  2703 => x"54",
  2704 => x"31",
  2705 => x"36",
  2706 => x"20",
  2707 => x"20",
  2708 => x"20",
  2709 => x"00",
  2710 => x"46",
  2711 => x"41",
  2712 => x"54",
  2713 => x"33",
  2714 => x"32",
  2715 => x"20",
  2716 => x"20",
  2717 => x"20",
  2718 => x"00",
  2719 => x"46",
  2720 => x"41",
  2721 => x"54",
  2722 => x"31",
  2723 => x"32",
  2724 => x"20",
  2725 => x"20",
  2726 => x"20",
  2727 => x"00",
  2728 => x"50",
  2729 => x"61",
  2730 => x"72",
  2731 => x"74",
  2732 => x"69",
  2733 => x"74",
  2734 => x"69",
  2735 => x"6f",
  2736 => x"6e",
  2737 => x"63",
  2738 => x"6f",
  2739 => x"75",
  2740 => x"6e",
  2741 => x"74",
  2742 => x"20",
  2743 => x"25",
  2744 => x"64",
  2745 => x"0a",
  2746 => x"00",
  2747 => x"48",
  2748 => x"75",
  2749 => x"6e",
  2750 => x"74",
  2751 => x"69",
  2752 => x"6e",
  2753 => x"67",
  2754 => x"20",
  2755 => x"66",
  2756 => x"6f",
  2757 => x"72",
  2758 => x"20",
  2759 => x"66",
  2760 => x"69",
  2761 => x"6c",
  2762 => x"65",
  2763 => x"73",
  2764 => x"79",
  2765 => x"73",
  2766 => x"74",
  2767 => x"65",
  2768 => x"6d",
  2769 => x"0a",
  2770 => x"00",
  2771 => x"46",
  2772 => x"41",
  2773 => x"54",
  2774 => x"33",
  2775 => x"32",
  2776 => x"20",
  2777 => x"20",
  2778 => x"20",
  2779 => x"00",
  2780 => x"46",
  2781 => x"41",
  2782 => x"54",
  2783 => x"31",
  2784 => x"36",
  2785 => x"20",
  2786 => x"20",
  2787 => x"20",
  2788 => x"00",
  2789 => x"52",
  2790 => x"65",
  2791 => x"61",
  2792 => x"64",
  2793 => x"69",
  2794 => x"6e",
  2795 => x"67",
  2796 => x"20",
  2797 => x"64",
  2798 => x"69",
  2799 => x"72",
  2800 => x"65",
  2801 => x"63",
  2802 => x"74",
  2803 => x"6f",
  2804 => x"72",
  2805 => x"79",
  2806 => x"20",
  2807 => x"73",
  2808 => x"65",
  2809 => x"63",
  2810 => x"74",
  2811 => x"6f",
  2812 => x"72",
  2813 => x"20",
  2814 => x"25",
  2815 => x"64",
  2816 => x"0a",
  2817 => x"00",
  2818 => x"66",
  2819 => x"69",
  2820 => x"6c",
  2821 => x"65",
  2822 => x"20",
  2823 => x"22",
  2824 => x"25",
  2825 => x"73",
  2826 => x"22",
  2827 => x"20",
  2828 => x"66",
  2829 => x"6f",
  2830 => x"75",
  2831 => x"6e",
  2832 => x"64",
  2833 => x"0d",
  2834 => x"00",
  2835 => x"47",
  2836 => x"65",
  2837 => x"74",
  2838 => x"46",
  2839 => x"41",
  2840 => x"54",
  2841 => x"4c",
  2842 => x"69",
  2843 => x"6e",
  2844 => x"6b",
  2845 => x"20",
  2846 => x"72",
  2847 => x"65",
  2848 => x"74",
  2849 => x"75",
  2850 => x"72",
  2851 => x"6e",
  2852 => x"65",
  2853 => x"64",
  2854 => x"20",
  2855 => x"25",
  2856 => x"64",
  2857 => x"0a",
  2858 => x"00",
  2859 => x"43",
  2860 => x"61",
  2861 => x"6e",
  2862 => x"27",
  2863 => x"74",
  2864 => x"20",
  2865 => x"6f",
  2866 => x"70",
  2867 => x"65",
  2868 => x"6e",
  2869 => x"20",
  2870 => x"25",
  2871 => x"73",
  2872 => x"0a",
  2873 => x"00",
  2874 => x"0e",
  2875 => x"5e",
  2876 => x"5b",
  2877 => x"5c",
  2878 => x"0e",
  2879 => x"c1",
  2880 => x"d0",
  2881 => x"fa",
  2882 => x"bf",
  2883 => x"02",
  2884 => x"ce",
  2885 => x"87",
  2886 => x"cc",
  2887 => x"66",
  2888 => x"4b",
  2889 => x"c7",
  2890 => x"b7",
  2891 => x"2b",
  2892 => x"cc",
  2893 => x"66",
  2894 => x"4c",
  2895 => x"c1",
  2896 => x"ff",
  2897 => x"9c",
  2898 => x"cc",
  2899 => x"87",
  2900 => x"cc",
  2901 => x"66",
  2902 => x"4b",
  2903 => x"c8",
  2904 => x"b7",
  2905 => x"2b",
  2906 => x"cc",
  2907 => x"66",
  2908 => x"4c",
  2909 => x"c3",
  2910 => x"ff",
  2911 => x"9c",
  2912 => x"c1",
  2913 => x"d1",
  2914 => x"ea",
  2915 => x"bf",
  2916 => x"ab",
  2917 => x"02",
  2918 => x"c0",
  2919 => x"e0",
  2920 => x"87",
  2921 => x"c1",
  2922 => x"c8",
  2923 => x"f2",
  2924 => x"1e",
  2925 => x"c1",
  2926 => x"d1",
  2927 => x"c6",
  2928 => x"bf",
  2929 => x"49",
  2930 => x"73",
  2931 => x"81",
  2932 => x"71",
  2933 => x"1e",
  2934 => x"e9",
  2935 => x"ef",
  2936 => x"87",
  2937 => x"c8",
  2938 => x"86",
  2939 => x"70",
  2940 => x"98",
  2941 => x"05",
  2942 => x"c5",
  2943 => x"87",
  2944 => x"c0",
  2945 => x"48",
  2946 => x"c0",
  2947 => x"fc",
  2948 => x"87",
  2949 => x"c1",
  2950 => x"d1",
  2951 => x"ee",
  2952 => x"5b",
  2953 => x"c1",
  2954 => x"d0",
  2955 => x"fa",
  2956 => x"bf",
  2957 => x"02",
  2958 => x"db",
  2959 => x"87",
  2960 => x"74",
  2961 => x"49",
  2962 => x"c4",
  2963 => x"91",
  2964 => x"c1",
  2965 => x"c8",
  2966 => x"f2",
  2967 => x"81",
  2968 => x"69",
  2969 => x"1e",
  2970 => x"eb",
  2971 => x"d5",
  2972 => x"87",
  2973 => x"c4",
  2974 => x"86",
  2975 => x"70",
  2976 => x"49",
  2977 => x"71",
  2978 => x"4a",
  2979 => x"cf",
  2980 => x"ff",
  2981 => x"ff",
  2982 => x"ff",
  2983 => x"ff",
  2984 => x"9a",
  2985 => x"d4",
  2986 => x"87",
  2987 => x"74",
  2988 => x"49",
  2989 => x"c2",
  2990 => x"91",
  2991 => x"c1",
  2992 => x"c8",
  2993 => x"f2",
  2994 => x"81",
  2995 => x"9f",
  2996 => x"69",
  2997 => x"49",
  2998 => x"71",
  2999 => x"1e",
  3000 => x"eb",
  3001 => x"e9",
  3002 => x"87",
  3003 => x"c4",
  3004 => x"86",
  3005 => x"70",
  3006 => x"4a",
  3007 => x"72",
  3008 => x"48",
  3009 => x"ec",
  3010 => x"fb",
  3011 => x"87",
  3012 => x"0e",
  3013 => x"5e",
  3014 => x"5b",
  3015 => x"5c",
  3016 => x"5d",
  3017 => x"0e",
  3018 => x"f8",
  3019 => x"86",
  3020 => x"c0",
  3021 => x"4b",
  3022 => x"c1",
  3023 => x"d1",
  3024 => x"ea",
  3025 => x"48",
  3026 => x"ff",
  3027 => x"78",
  3028 => x"c1",
  3029 => x"d1",
  3030 => x"ce",
  3031 => x"bf",
  3032 => x"4d",
  3033 => x"c1",
  3034 => x"d1",
  3035 => x"d2",
  3036 => x"bf",
  3037 => x"4c",
  3038 => x"c1",
  3039 => x"d0",
  3040 => x"fa",
  3041 => x"bf",
  3042 => x"02",
  3043 => x"c9",
  3044 => x"87",
  3045 => x"c1",
  3046 => x"d0",
  3047 => x"f2",
  3048 => x"bf",
  3049 => x"49",
  3050 => x"c4",
  3051 => x"31",
  3052 => x"c7",
  3053 => x"87",
  3054 => x"c1",
  3055 => x"d1",
  3056 => x"d6",
  3057 => x"bf",
  3058 => x"49",
  3059 => x"c4",
  3060 => x"31",
  3061 => x"c4",
  3062 => x"a6",
  3063 => x"59",
  3064 => x"c4",
  3065 => x"a6",
  3066 => x"48",
  3067 => x"c0",
  3068 => x"78",
  3069 => x"6e",
  3070 => x"48",
  3071 => x"c0",
  3072 => x"a8",
  3073 => x"06",
  3074 => x"c3",
  3075 => x"d5",
  3076 => x"87",
  3077 => x"c4",
  3078 => x"66",
  3079 => x"49",
  3080 => x"cf",
  3081 => x"99",
  3082 => x"05",
  3083 => x"dc",
  3084 => x"87",
  3085 => x"74",
  3086 => x"1e",
  3087 => x"c0",
  3088 => x"eb",
  3089 => x"e5",
  3090 => x"1e",
  3091 => x"d5",
  3092 => x"f7",
  3093 => x"87",
  3094 => x"c1",
  3095 => x"c8",
  3096 => x"f2",
  3097 => x"1e",
  3098 => x"74",
  3099 => x"1e",
  3100 => x"c1",
  3101 => x"84",
  3102 => x"e7",
  3103 => x"c7",
  3104 => x"87",
  3105 => x"d0",
  3106 => x"86",
  3107 => x"c1",
  3108 => x"c8",
  3109 => x"f2",
  3110 => x"4b",
  3111 => x"c3",
  3112 => x"87",
  3113 => x"c0",
  3114 => x"e0",
  3115 => x"83",
  3116 => x"97",
  3117 => x"6b",
  3118 => x"49",
  3119 => x"71",
  3120 => x"99",
  3121 => x"02",
  3122 => x"c2",
  3123 => x"d4",
  3124 => x"87",
  3125 => x"97",
  3126 => x"6b",
  3127 => x"49",
  3128 => x"c3",
  3129 => x"e5",
  3130 => x"a9",
  3131 => x"02",
  3132 => x"c2",
  3133 => x"ca",
  3134 => x"87",
  3135 => x"cb",
  3136 => x"a3",
  3137 => x"49",
  3138 => x"97",
  3139 => x"69",
  3140 => x"49",
  3141 => x"d8",
  3142 => x"99",
  3143 => x"05",
  3144 => x"c1",
  3145 => x"fe",
  3146 => x"87",
  3147 => x"cb",
  3148 => x"1e",
  3149 => x"c0",
  3150 => x"e0",
  3151 => x"66",
  3152 => x"1e",
  3153 => x"73",
  3154 => x"1e",
  3155 => x"e9",
  3156 => x"e6",
  3157 => x"87",
  3158 => x"cc",
  3159 => x"86",
  3160 => x"70",
  3161 => x"98",
  3162 => x"05",
  3163 => x"c1",
  3164 => x"eb",
  3165 => x"87",
  3166 => x"dc",
  3167 => x"a3",
  3168 => x"49",
  3169 => x"69",
  3170 => x"1e",
  3171 => x"e8",
  3172 => x"cc",
  3173 => x"87",
  3174 => x"70",
  3175 => x"4a",
  3176 => x"dc",
  3177 => x"66",
  3178 => x"49",
  3179 => x"c4",
  3180 => x"81",
  3181 => x"72",
  3182 => x"79",
  3183 => x"da",
  3184 => x"a3",
  3185 => x"49",
  3186 => x"9f",
  3187 => x"69",
  3188 => x"49",
  3189 => x"71",
  3190 => x"1e",
  3191 => x"e8",
  3192 => x"ea",
  3193 => x"87",
  3194 => x"c8",
  3195 => x"86",
  3196 => x"c4",
  3197 => x"a6",
  3198 => x"58",
  3199 => x"c1",
  3200 => x"d0",
  3201 => x"fa",
  3202 => x"bf",
  3203 => x"02",
  3204 => x"dc",
  3205 => x"87",
  3206 => x"d4",
  3207 => x"a3",
  3208 => x"49",
  3209 => x"9f",
  3210 => x"69",
  3211 => x"49",
  3212 => x"71",
  3213 => x"1e",
  3214 => x"e8",
  3215 => x"d3",
  3216 => x"87",
  3217 => x"c4",
  3218 => x"86",
  3219 => x"70",
  3220 => x"49",
  3221 => x"c0",
  3222 => x"ff",
  3223 => x"ff",
  3224 => x"99",
  3225 => x"71",
  3226 => x"48",
  3227 => x"d0",
  3228 => x"30",
  3229 => x"c8",
  3230 => x"a6",
  3231 => x"58",
  3232 => x"c5",
  3233 => x"87",
  3234 => x"c4",
  3235 => x"a6",
  3236 => x"48",
  3237 => x"c0",
  3238 => x"78",
  3239 => x"c4",
  3240 => x"66",
  3241 => x"4a",
  3242 => x"6e",
  3243 => x"82",
  3244 => x"d8",
  3245 => x"66",
  3246 => x"49",
  3247 => x"c8",
  3248 => x"81",
  3249 => x"72",
  3250 => x"79",
  3251 => x"d8",
  3252 => x"66",
  3253 => x"48",
  3254 => x"c0",
  3255 => x"78",
  3256 => x"dc",
  3257 => x"66",
  3258 => x"1e",
  3259 => x"c0",
  3260 => x"ec",
  3261 => x"c2",
  3262 => x"1e",
  3263 => x"d3",
  3264 => x"cb",
  3265 => x"87",
  3266 => x"c8",
  3267 => x"86",
  3268 => x"c1",
  3269 => x"48",
  3270 => x"c1",
  3271 => x"cc",
  3272 => x"87",
  3273 => x"c4",
  3274 => x"66",
  3275 => x"48",
  3276 => x"c1",
  3277 => x"80",
  3278 => x"c8",
  3279 => x"a6",
  3280 => x"58",
  3281 => x"c4",
  3282 => x"66",
  3283 => x"48",
  3284 => x"6e",
  3285 => x"a8",
  3286 => x"04",
  3287 => x"fc",
  3288 => x"eb",
  3289 => x"87",
  3290 => x"c1",
  3291 => x"d0",
  3292 => x"fa",
  3293 => x"bf",
  3294 => x"02",
  3295 => x"c0",
  3296 => x"f1",
  3297 => x"87",
  3298 => x"75",
  3299 => x"1e",
  3300 => x"f9",
  3301 => x"d3",
  3302 => x"87",
  3303 => x"70",
  3304 => x"4d",
  3305 => x"75",
  3306 => x"1e",
  3307 => x"c0",
  3308 => x"ec",
  3309 => x"d3",
  3310 => x"1e",
  3311 => x"d2",
  3312 => x"db",
  3313 => x"87",
  3314 => x"cc",
  3315 => x"86",
  3316 => x"75",
  3317 => x"49",
  3318 => x"cf",
  3319 => x"ff",
  3320 => x"ff",
  3321 => x"ff",
  3322 => x"f8",
  3323 => x"99",
  3324 => x"a9",
  3325 => x"02",
  3326 => x"d3",
  3327 => x"87",
  3328 => x"75",
  3329 => x"49",
  3330 => x"c2",
  3331 => x"89",
  3332 => x"c1",
  3333 => x"d0",
  3334 => x"f2",
  3335 => x"bf",
  3336 => x"91",
  3337 => x"c1",
  3338 => x"d1",
  3339 => x"ca",
  3340 => x"bf",
  3341 => x"4c",
  3342 => x"71",
  3343 => x"84",
  3344 => x"fb",
  3345 => x"e5",
  3346 => x"87",
  3347 => x"c0",
  3348 => x"48",
  3349 => x"f8",
  3350 => x"8e",
  3351 => x"e7",
  3352 => x"e3",
  3353 => x"87",
  3354 => x"0e",
  3355 => x"5e",
  3356 => x"5b",
  3357 => x"5c",
  3358 => x"5d",
  3359 => x"0e",
  3360 => x"d0",
  3361 => x"66",
  3362 => x"1e",
  3363 => x"c1",
  3364 => x"d1",
  3365 => x"ee",
  3366 => x"1e",
  3367 => x"fa",
  3368 => x"da",
  3369 => x"87",
  3370 => x"c8",
  3371 => x"86",
  3372 => x"70",
  3373 => x"98",
  3374 => x"02",
  3375 => x"c1",
  3376 => x"f5",
  3377 => x"87",
  3378 => x"c1",
  3379 => x"d1",
  3380 => x"f2",
  3381 => x"bf",
  3382 => x"49",
  3383 => x"c7",
  3384 => x"ff",
  3385 => x"81",
  3386 => x"c9",
  3387 => x"29",
  3388 => x"71",
  3389 => x"4d",
  3390 => x"c0",
  3391 => x"4c",
  3392 => x"4b",
  3393 => x"b7",
  3394 => x"ad",
  3395 => x"06",
  3396 => x"c1",
  3397 => x"f0",
  3398 => x"87",
  3399 => x"c1",
  3400 => x"d1",
  3401 => x"ca",
  3402 => x"bf",
  3403 => x"49",
  3404 => x"c1",
  3405 => x"d1",
  3406 => x"f6",
  3407 => x"bf",
  3408 => x"4a",
  3409 => x"c2",
  3410 => x"8a",
  3411 => x"c1",
  3412 => x"d0",
  3413 => x"f2",
  3414 => x"bf",
  3415 => x"92",
  3416 => x"72",
  3417 => x"a1",
  3418 => x"49",
  3419 => x"c1",
  3420 => x"d0",
  3421 => x"f6",
  3422 => x"bf",
  3423 => x"4a",
  3424 => x"73",
  3425 => x"9a",
  3426 => x"72",
  3427 => x"a1",
  3428 => x"49",
  3429 => x"d4",
  3430 => x"66",
  3431 => x"1e",
  3432 => x"71",
  3433 => x"1e",
  3434 => x"e1",
  3435 => x"fb",
  3436 => x"87",
  3437 => x"c8",
  3438 => x"86",
  3439 => x"70",
  3440 => x"98",
  3441 => x"05",
  3442 => x"c5",
  3443 => x"87",
  3444 => x"c0",
  3445 => x"48",
  3446 => x"c1",
  3447 => x"c3",
  3448 => x"87",
  3449 => x"c1",
  3450 => x"83",
  3451 => x"c1",
  3452 => x"d0",
  3453 => x"f6",
  3454 => x"bf",
  3455 => x"49",
  3456 => x"73",
  3457 => x"99",
  3458 => x"05",
  3459 => x"ce",
  3460 => x"87",
  3461 => x"c1",
  3462 => x"d1",
  3463 => x"f6",
  3464 => x"bf",
  3465 => x"1e",
  3466 => x"f6",
  3467 => x"ed",
  3468 => x"87",
  3469 => x"c4",
  3470 => x"86",
  3471 => x"c1",
  3472 => x"d1",
  3473 => x"fa",
  3474 => x"58",
  3475 => x"d4",
  3476 => x"66",
  3477 => x"48",
  3478 => x"c8",
  3479 => x"c0",
  3480 => x"80",
  3481 => x"d8",
  3482 => x"a6",
  3483 => x"58",
  3484 => x"c1",
  3485 => x"84",
  3486 => x"75",
  3487 => x"b7",
  3488 => x"ac",
  3489 => x"04",
  3490 => x"fe",
  3491 => x"e2",
  3492 => x"87",
  3493 => x"d0",
  3494 => x"87",
  3495 => x"d0",
  3496 => x"66",
  3497 => x"1e",
  3498 => x"c0",
  3499 => x"ec",
  3500 => x"eb",
  3501 => x"1e",
  3502 => x"cf",
  3503 => x"dc",
  3504 => x"87",
  3505 => x"c8",
  3506 => x"86",
  3507 => x"c0",
  3508 => x"48",
  3509 => x"c5",
  3510 => x"87",
  3511 => x"c1",
  3512 => x"d1",
  3513 => x"f2",
  3514 => x"bf",
  3515 => x"48",
  3516 => x"e4",
  3517 => x"fe",
  3518 => x"87",
  3519 => x"1e",
  3520 => x"c0",
  3521 => x"f6",
  3522 => x"e8",
  3523 => x"c0",
  3524 => x"c0",
  3525 => x"48",
  3526 => x"c4",
  3527 => x"66",
  3528 => x"50",
  3529 => x"48",
  3530 => x"26",
  3531 => x"4f",
  3532 => x"0e",
  3533 => x"5e",
  3534 => x"5b",
  3535 => x"5c",
  3536 => x"0e",
  3537 => x"cc",
  3538 => x"66",
  3539 => x"4c",
  3540 => x"c0",
  3541 => x"4b",
  3542 => x"14",
  3543 => x"49",
  3544 => x"71",
  3545 => x"99",
  3546 => x"02",
  3547 => x"d0",
  3548 => x"87",
  3549 => x"71",
  3550 => x"1e",
  3551 => x"ff",
  3552 => x"dd",
  3553 => x"87",
  3554 => x"c4",
  3555 => x"86",
  3556 => x"c1",
  3557 => x"83",
  3558 => x"14",
  3559 => x"49",
  3560 => x"71",
  3561 => x"99",
  3562 => x"05",
  3563 => x"f0",
  3564 => x"87",
  3565 => x"73",
  3566 => x"48",
  3567 => x"c2",
  3568 => x"87",
  3569 => x"26",
  3570 => x"4d",
  3571 => x"26",
  3572 => x"4c",
  3573 => x"26",
  3574 => x"4b",
  3575 => x"26",
  3576 => x"4f",
  3577 => x"0e",
  3578 => x"5e",
  3579 => x"5b",
  3580 => x"5c",
  3581 => x"5d",
  3582 => x"0e",
  3583 => x"1e",
  3584 => x"d8",
  3585 => x"66",
  3586 => x"4b",
  3587 => x"d4",
  3588 => x"66",
  3589 => x"4a",
  3590 => x"c0",
  3591 => x"4c",
  3592 => x"b7",
  3593 => x"ab",
  3594 => x"06",
  3595 => x"c1",
  3596 => x"ca",
  3597 => x"87",
  3598 => x"12",
  3599 => x"49",
  3600 => x"c8",
  3601 => x"31",
  3602 => x"c1",
  3603 => x"8b",
  3604 => x"c0",
  3605 => x"b7",
  3606 => x"ab",
  3607 => x"06",
  3608 => x"c7",
  3609 => x"87",
  3610 => x"12",
  3611 => x"48",
  3612 => x"c4",
  3613 => x"a6",
  3614 => x"58",
  3615 => x"c2",
  3616 => x"87",
  3617 => x"c0",
  3618 => x"7e",
  3619 => x"6e",
  3620 => x"b1",
  3621 => x"c8",
  3622 => x"31",
  3623 => x"c1",
  3624 => x"8b",
  3625 => x"c0",
  3626 => x"b7",
  3627 => x"ab",
  3628 => x"06",
  3629 => x"c4",
  3630 => x"87",
  3631 => x"12",
  3632 => x"4d",
  3633 => x"c2",
  3634 => x"87",
  3635 => x"c0",
  3636 => x"4d",
  3637 => x"75",
  3638 => x"b1",
  3639 => x"c8",
  3640 => x"31",
  3641 => x"c1",
  3642 => x"8b",
  3643 => x"c0",
  3644 => x"b7",
  3645 => x"ab",
  3646 => x"06",
  3647 => x"c7",
  3648 => x"87",
  3649 => x"12",
  3650 => x"48",
  3651 => x"c4",
  3652 => x"a6",
  3653 => x"58",
  3654 => x"c2",
  3655 => x"87",
  3656 => x"c0",
  3657 => x"7e",
  3658 => x"6e",
  3659 => x"b1",
  3660 => x"71",
  3661 => x"a4",
  3662 => x"4c",
  3663 => x"c1",
  3664 => x"8b",
  3665 => x"c0",
  3666 => x"b7",
  3667 => x"ab",
  3668 => x"01",
  3669 => x"fe",
  3670 => x"f6",
  3671 => x"87",
  3672 => x"74",
  3673 => x"48",
  3674 => x"26",
  3675 => x"26",
  3676 => x"4d",
  3677 => x"26",
  3678 => x"4c",
  3679 => x"26",
  3680 => x"4b",
  3681 => x"26",
  3682 => x"4f",
  3683 => x"0e",
  3684 => x"5e",
  3685 => x"5b",
  3686 => x"5c",
  3687 => x"5d",
  3688 => x"0e",
  3689 => x"1e",
  3690 => x"d8",
  3691 => x"66",
  3692 => x"4c",
  3693 => x"d4",
  3694 => x"66",
  3695 => x"4b",
  3696 => x"c2",
  3697 => x"2c",
  3698 => x"74",
  3699 => x"49",
  3700 => x"c1",
  3701 => x"8c",
  3702 => x"71",
  3703 => x"99",
  3704 => x"02",
  3705 => x"c1",
  3706 => x"ca",
  3707 => x"87",
  3708 => x"23",
  3709 => x"7e",
  3710 => x"c0",
  3711 => x"4d",
  3712 => x"6e",
  3713 => x"49",
  3714 => x"dc",
  3715 => x"29",
  3716 => x"c0",
  3717 => x"f0",
  3718 => x"81",
  3719 => x"c0",
  3720 => x"f9",
  3721 => x"a9",
  3722 => x"06",
  3723 => x"c2",
  3724 => x"87",
  3725 => x"c7",
  3726 => x"81",
  3727 => x"71",
  3728 => x"1e",
  3729 => x"fc",
  3730 => x"eb",
  3731 => x"87",
  3732 => x"c4",
  3733 => x"86",
  3734 => x"6e",
  3735 => x"48",
  3736 => x"c4",
  3737 => x"30",
  3738 => x"c4",
  3739 => x"a6",
  3740 => x"58",
  3741 => x"c1",
  3742 => x"85",
  3743 => x"c8",
  3744 => x"b7",
  3745 => x"ad",
  3746 => x"04",
  3747 => x"ff",
  3748 => x"da",
  3749 => x"87",
  3750 => x"c0",
  3751 => x"e0",
  3752 => x"1e",
  3753 => x"fc",
  3754 => x"d3",
  3755 => x"87",
  3756 => x"c4",
  3757 => x"86",
  3758 => x"74",
  3759 => x"49",
  3760 => x"c3",
  3761 => x"99",
  3762 => x"05",
  3763 => x"c7",
  3764 => x"87",
  3765 => x"ca",
  3766 => x"1e",
  3767 => x"fc",
  3768 => x"c5",
  3769 => x"87",
  3770 => x"c4",
  3771 => x"86",
  3772 => x"74",
  3773 => x"49",
  3774 => x"c1",
  3775 => x"8c",
  3776 => x"71",
  3777 => x"99",
  3778 => x"05",
  3779 => x"fe",
  3780 => x"f6",
  3781 => x"87",
  3782 => x"ca",
  3783 => x"1e",
  3784 => x"fb",
  3785 => x"f4",
  3786 => x"87",
  3787 => x"f8",
  3788 => x"8e",
  3789 => x"26",
  3790 => x"4d",
  3791 => x"26",
  3792 => x"4c",
  3793 => x"26",
  3794 => x"4b",
  3795 => x"26",
  3796 => x"4f",
  3797 => x"0e",
  3798 => x"5e",
  3799 => x"5b",
  3800 => x"5c",
  3801 => x"5d",
  3802 => x"0e",
  3803 => x"d0",
  3804 => x"66",
  3805 => x"4c",
  3806 => x"c0",
  3807 => x"e0",
  3808 => x"66",
  3809 => x"4a",
  3810 => x"c1",
  3811 => x"d1",
  3812 => x"fa",
  3813 => x"4b",
  3814 => x"c0",
  3815 => x"4d",
  3816 => x"74",
  3817 => x"9c",
  3818 => x"05",
  3819 => x"ce",
  3820 => x"87",
  3821 => x"c1",
  3822 => x"d1",
  3823 => x"fb",
  3824 => x"4b",
  3825 => x"c1",
  3826 => x"d1",
  3827 => x"fa",
  3828 => x"48",
  3829 => x"c0",
  3830 => x"f0",
  3831 => x"50",
  3832 => x"c1",
  3833 => x"d5",
  3834 => x"87",
  3835 => x"74",
  3836 => x"9c",
  3837 => x"02",
  3838 => x"c0",
  3839 => x"ec",
  3840 => x"87",
  3841 => x"72",
  3842 => x"1e",
  3843 => x"74",
  3844 => x"49",
  3845 => x"d8",
  3846 => x"66",
  3847 => x"4a",
  3848 => x"ca",
  3849 => x"d6",
  3850 => x"87",
  3851 => x"26",
  3852 => x"4a",
  3853 => x"c0",
  3854 => x"fd",
  3855 => x"fc",
  3856 => x"81",
  3857 => x"11",
  3858 => x"53",
  3859 => x"71",
  3860 => x"1e",
  3861 => x"72",
  3862 => x"1e",
  3863 => x"74",
  3864 => x"49",
  3865 => x"dc",
  3866 => x"66",
  3867 => x"4a",
  3868 => x"ca",
  3869 => x"c2",
  3870 => x"87",
  3871 => x"70",
  3872 => x"4c",
  3873 => x"26",
  3874 => x"4a",
  3875 => x"26",
  3876 => x"49",
  3877 => x"c1",
  3878 => x"8a",
  3879 => x"74",
  3880 => x"9c",
  3881 => x"05",
  3882 => x"ff",
  3883 => x"d4",
  3884 => x"87",
  3885 => x"c0",
  3886 => x"b7",
  3887 => x"aa",
  3888 => x"06",
  3889 => x"dd",
  3890 => x"87",
  3891 => x"c0",
  3892 => x"e4",
  3893 => x"66",
  3894 => x"02",
  3895 => x"c5",
  3896 => x"87",
  3897 => x"c0",
  3898 => x"f0",
  3899 => x"49",
  3900 => x"c3",
  3901 => x"87",
  3902 => x"c0",
  3903 => x"e0",
  3904 => x"49",
  3905 => x"73",
  3906 => x"09",
  3907 => x"97",
  3908 => x"79",
  3909 => x"09",
  3910 => x"c1",
  3911 => x"83",
  3912 => x"8a",
  3913 => x"c0",
  3914 => x"b7",
  3915 => x"aa",
  3916 => x"01",
  3917 => x"ff",
  3918 => x"e3",
  3919 => x"87",
  3920 => x"c1",
  3921 => x"d1",
  3922 => x"fa",
  3923 => x"ab",
  3924 => x"02",
  3925 => x"db",
  3926 => x"87",
  3927 => x"d8",
  3928 => x"66",
  3929 => x"4c",
  3930 => x"dc",
  3931 => x"66",
  3932 => x"1e",
  3933 => x"c1",
  3934 => x"8b",
  3935 => x"97",
  3936 => x"6b",
  3937 => x"49",
  3938 => x"71",
  3939 => x"1e",
  3940 => x"74",
  3941 => x"0f",
  3942 => x"c8",
  3943 => x"86",
  3944 => x"c1",
  3945 => x"85",
  3946 => x"c1",
  3947 => x"d1",
  3948 => x"fa",
  3949 => x"ab",
  3950 => x"05",
  3951 => x"ff",
  3952 => x"e8",
  3953 => x"87",
  3954 => x"75",
  3955 => x"48",
  3956 => x"26",
  3957 => x"4d",
  3958 => x"26",
  3959 => x"4c",
  3960 => x"26",
  3961 => x"4b",
  3962 => x"26",
  3963 => x"4f",
  3964 => x"30",
  3965 => x"31",
  3966 => x"32",
  3967 => x"33",
  3968 => x"34",
  3969 => x"35",
  3970 => x"36",
  3971 => x"37",
  3972 => x"38",
  3973 => x"39",
  3974 => x"41",
  3975 => x"42",
  3976 => x"43",
  3977 => x"44",
  3978 => x"45",
  3979 => x"46",
  3980 => x"00",
  3981 => x"0e",
  3982 => x"5e",
  3983 => x"5b",
  3984 => x"5c",
  3985 => x"5d",
  3986 => x"0e",
  3987 => x"d0",
  3988 => x"66",
  3989 => x"4c",
  3990 => x"ff",
  3991 => x"4d",
  3992 => x"14",
  3993 => x"4b",
  3994 => x"73",
  3995 => x"9b",
  3996 => x"02",
  3997 => x"d8",
  3998 => x"87",
  3999 => x"c1",
  4000 => x"85",
  4001 => x"d8",
  4002 => x"66",
  4003 => x"1e",
  4004 => x"73",
  4005 => x"1e",
  4006 => x"dc",
  4007 => x"66",
  4008 => x"0f",
  4009 => x"c8",
  4010 => x"86",
  4011 => x"73",
  4012 => x"a8",
  4013 => x"05",
  4014 => x"c7",
  4015 => x"87",
  4016 => x"14",
  4017 => x"4b",
  4018 => x"73",
  4019 => x"9b",
  4020 => x"05",
  4021 => x"e8",
  4022 => x"87",
  4023 => x"75",
  4024 => x"48",
  4025 => x"26",
  4026 => x"4d",
  4027 => x"26",
  4028 => x"4c",
  4029 => x"26",
  4030 => x"4b",
  4031 => x"26",
  4032 => x"4f",
  4033 => x"0e",
  4034 => x"5e",
  4035 => x"5b",
  4036 => x"5c",
  4037 => x"5d",
  4038 => x"0e",
  4039 => x"ec",
  4040 => x"86",
  4041 => x"c0",
  4042 => x"e8",
  4043 => x"66",
  4044 => x"4d",
  4045 => x"c0",
  4046 => x"4c",
  4047 => x"c4",
  4048 => x"a6",
  4049 => x"48",
  4050 => x"c0",
  4051 => x"78",
  4052 => x"c0",
  4053 => x"e4",
  4054 => x"66",
  4055 => x"97",
  4056 => x"bf",
  4057 => x"4b",
  4058 => x"c0",
  4059 => x"e4",
  4060 => x"66",
  4061 => x"48",
  4062 => x"c1",
  4063 => x"80",
  4064 => x"c0",
  4065 => x"e8",
  4066 => x"a6",
  4067 => x"58",
  4068 => x"73",
  4069 => x"9b",
  4070 => x"02",
  4071 => x"c6",
  4072 => x"d7",
  4073 => x"87",
  4074 => x"c4",
  4075 => x"66",
  4076 => x"02",
  4077 => x"c5",
  4078 => x"d9",
  4079 => x"87",
  4080 => x"c8",
  4081 => x"a6",
  4082 => x"48",
  4083 => x"c0",
  4084 => x"78",
  4085 => x"fc",
  4086 => x"80",
  4087 => x"c0",
  4088 => x"78",
  4089 => x"73",
  4090 => x"49",
  4091 => x"c0",
  4092 => x"e0",
  4093 => x"89",
  4094 => x"02",
  4095 => x"c3",
  4096 => x"c6",
  4097 => x"87",
  4098 => x"c3",
  4099 => x"89",
  4100 => x"02",
  4101 => x"c3",
  4102 => x"c0",
  4103 => x"87",
  4104 => x"c2",
  4105 => x"89",
  4106 => x"02",
  4107 => x"c2",
  4108 => x"e8",
  4109 => x"87",
  4110 => x"c2",
  4111 => x"89",
  4112 => x"02",
  4113 => x"c2",
  4114 => x"f4",
  4115 => x"87",
  4116 => x"c4",
  4117 => x"89",
  4118 => x"02",
  4119 => x"c2",
  4120 => x"ee",
  4121 => x"87",
  4122 => x"c2",
  4123 => x"89",
  4124 => x"02",
  4125 => x"c2",
  4126 => x"e8",
  4127 => x"87",
  4128 => x"c3",
  4129 => x"89",
  4130 => x"02",
  4131 => x"c2",
  4132 => x"ea",
  4133 => x"87",
  4134 => x"d4",
  4135 => x"89",
  4136 => x"02",
  4137 => x"c0",
  4138 => x"f6",
  4139 => x"87",
  4140 => x"d4",
  4141 => x"89",
  4142 => x"02",
  4143 => x"c1",
  4144 => x"c0",
  4145 => x"87",
  4146 => x"ca",
  4147 => x"89",
  4148 => x"02",
  4149 => x"c0",
  4150 => x"f2",
  4151 => x"87",
  4152 => x"c1",
  4153 => x"89",
  4154 => x"02",
  4155 => x"c1",
  4156 => x"e1",
  4157 => x"87",
  4158 => x"c1",
  4159 => x"89",
  4160 => x"02",
  4161 => x"df",
  4162 => x"87",
  4163 => x"c8",
  4164 => x"89",
  4165 => x"02",
  4166 => x"c1",
  4167 => x"ce",
  4168 => x"87",
  4169 => x"c4",
  4170 => x"89",
  4171 => x"02",
  4172 => x"c0",
  4173 => x"e3",
  4174 => x"87",
  4175 => x"c3",
  4176 => x"89",
  4177 => x"02",
  4178 => x"c0",
  4179 => x"e5",
  4180 => x"87",
  4181 => x"c2",
  4182 => x"89",
  4183 => x"02",
  4184 => x"c8",
  4185 => x"87",
  4186 => x"c3",
  4187 => x"89",
  4188 => x"02",
  4189 => x"d3",
  4190 => x"87",
  4191 => x"c1",
  4192 => x"fa",
  4193 => x"87",
  4194 => x"c8",
  4195 => x"a6",
  4196 => x"48",
  4197 => x"ca",
  4198 => x"78",
  4199 => x"c2",
  4200 => x"d2",
  4201 => x"87",
  4202 => x"c8",
  4203 => x"a6",
  4204 => x"48",
  4205 => x"c2",
  4206 => x"78",
  4207 => x"c2",
  4208 => x"ca",
  4209 => x"87",
  4210 => x"c8",
  4211 => x"a6",
  4212 => x"48",
  4213 => x"d0",
  4214 => x"78",
  4215 => x"c2",
  4216 => x"c2",
  4217 => x"87",
  4218 => x"c0",
  4219 => x"f0",
  4220 => x"66",
  4221 => x"1e",
  4222 => x"c0",
  4223 => x"f0",
  4224 => x"66",
  4225 => x"1e",
  4226 => x"c4",
  4227 => x"85",
  4228 => x"75",
  4229 => x"49",
  4230 => x"c4",
  4231 => x"89",
  4232 => x"69",
  4233 => x"1e",
  4234 => x"fc",
  4235 => x"c0",
  4236 => x"87",
  4237 => x"cc",
  4238 => x"86",
  4239 => x"70",
  4240 => x"49",
  4241 => x"71",
  4242 => x"a4",
  4243 => x"4c",
  4244 => x"c1",
  4245 => x"e5",
  4246 => x"87",
  4247 => x"c4",
  4248 => x"a6",
  4249 => x"48",
  4250 => x"c1",
  4251 => x"78",
  4252 => x"c1",
  4253 => x"dd",
  4254 => x"87",
  4255 => x"c0",
  4256 => x"f0",
  4257 => x"66",
  4258 => x"1e",
  4259 => x"c4",
  4260 => x"85",
  4261 => x"75",
  4262 => x"49",
  4263 => x"c4",
  4264 => x"89",
  4265 => x"69",
  4266 => x"1e",
  4267 => x"c0",
  4268 => x"f4",
  4269 => x"66",
  4270 => x"0f",
  4271 => x"c8",
  4272 => x"86",
  4273 => x"c1",
  4274 => x"84",
  4275 => x"c1",
  4276 => x"c6",
  4277 => x"87",
  4278 => x"c0",
  4279 => x"f0",
  4280 => x"66",
  4281 => x"1e",
  4282 => x"c0",
  4283 => x"e5",
  4284 => x"1e",
  4285 => x"c0",
  4286 => x"f4",
  4287 => x"66",
  4288 => x"0f",
  4289 => x"c8",
  4290 => x"86",
  4291 => x"c1",
  4292 => x"84",
  4293 => x"c0",
  4294 => x"f4",
  4295 => x"87",
  4296 => x"c4",
  4297 => x"a6",
  4298 => x"48",
  4299 => x"c1",
  4300 => x"78",
  4301 => x"c0",
  4302 => x"ec",
  4303 => x"87",
  4304 => x"cc",
  4305 => x"a6",
  4306 => x"48",
  4307 => x"c1",
  4308 => x"78",
  4309 => x"f8",
  4310 => x"80",
  4311 => x"c1",
  4312 => x"78",
  4313 => x"c0",
  4314 => x"e0",
  4315 => x"87",
  4316 => x"c0",
  4317 => x"f0",
  4318 => x"ab",
  4319 => x"06",
  4320 => x"da",
  4321 => x"87",
  4322 => x"c0",
  4323 => x"f9",
  4324 => x"ab",
  4325 => x"03",
  4326 => x"d4",
  4327 => x"87",
  4328 => x"d0",
  4329 => x"66",
  4330 => x"49",
  4331 => x"ca",
  4332 => x"91",
  4333 => x"73",
  4334 => x"4a",
  4335 => x"c0",
  4336 => x"f0",
  4337 => x"8a",
  4338 => x"d0",
  4339 => x"a6",
  4340 => x"48",
  4341 => x"72",
  4342 => x"a1",
  4343 => x"78",
  4344 => x"f4",
  4345 => x"80",
  4346 => x"c1",
  4347 => x"78",
  4348 => x"c8",
  4349 => x"66",
  4350 => x"02",
  4351 => x"c1",
  4352 => x"e9",
  4353 => x"87",
  4354 => x"c4",
  4355 => x"85",
  4356 => x"75",
  4357 => x"49",
  4358 => x"c4",
  4359 => x"89",
  4360 => x"69",
  4361 => x"7e",
  4362 => x"c1",
  4363 => x"e4",
  4364 => x"ab",
  4365 => x"05",
  4366 => x"d8",
  4367 => x"87",
  4368 => x"6e",
  4369 => x"48",
  4370 => x"c0",
  4371 => x"b7",
  4372 => x"a8",
  4373 => x"03",
  4374 => x"d0",
  4375 => x"87",
  4376 => x"c0",
  4377 => x"ed",
  4378 => x"1e",
  4379 => x"f2",
  4380 => x"e1",
  4381 => x"87",
  4382 => x"c4",
  4383 => x"86",
  4384 => x"6e",
  4385 => x"48",
  4386 => x"c0",
  4387 => x"08",
  4388 => x"88",
  4389 => x"c4",
  4390 => x"a6",
  4391 => x"58",
  4392 => x"cc",
  4393 => x"66",
  4394 => x"1e",
  4395 => x"d4",
  4396 => x"66",
  4397 => x"1e",
  4398 => x"c0",
  4399 => x"f8",
  4400 => x"66",
  4401 => x"1e",
  4402 => x"c0",
  4403 => x"f8",
  4404 => x"66",
  4405 => x"1e",
  4406 => x"d8",
  4407 => x"66",
  4408 => x"1e",
  4409 => x"d4",
  4410 => x"66",
  4411 => x"1e",
  4412 => x"f6",
  4413 => x"d6",
  4414 => x"87",
  4415 => x"d8",
  4416 => x"86",
  4417 => x"70",
  4418 => x"49",
  4419 => x"71",
  4420 => x"a4",
  4421 => x"4c",
  4422 => x"c0",
  4423 => x"e2",
  4424 => x"87",
  4425 => x"c0",
  4426 => x"e5",
  4427 => x"ab",
  4428 => x"05",
  4429 => x"d0",
  4430 => x"87",
  4431 => x"cc",
  4432 => x"a6",
  4433 => x"48",
  4434 => x"c0",
  4435 => x"78",
  4436 => x"c4",
  4437 => x"80",
  4438 => x"c0",
  4439 => x"78",
  4440 => x"c4",
  4441 => x"a6",
  4442 => x"48",
  4443 => x"c1",
  4444 => x"78",
  4445 => x"cc",
  4446 => x"87",
  4447 => x"c0",
  4448 => x"f0",
  4449 => x"66",
  4450 => x"1e",
  4451 => x"73",
  4452 => x"1e",
  4453 => x"c0",
  4454 => x"f4",
  4455 => x"66",
  4456 => x"0f",
  4457 => x"c8",
  4458 => x"86",
  4459 => x"c0",
  4460 => x"e4",
  4461 => x"66",
  4462 => x"97",
  4463 => x"bf",
  4464 => x"4b",
  4465 => x"c0",
  4466 => x"e4",
  4467 => x"66",
  4468 => x"48",
  4469 => x"c1",
  4470 => x"80",
  4471 => x"c0",
  4472 => x"e8",
  4473 => x"a6",
  4474 => x"58",
  4475 => x"73",
  4476 => x"9b",
  4477 => x"05",
  4478 => x"f9",
  4479 => x"e9",
  4480 => x"87",
  4481 => x"74",
  4482 => x"48",
  4483 => x"ec",
  4484 => x"8e",
  4485 => x"26",
  4486 => x"4d",
  4487 => x"26",
  4488 => x"4c",
  4489 => x"26",
  4490 => x"4b",
  4491 => x"26",
  4492 => x"4f",
  4493 => x"1e",
  4494 => x"c0",
  4495 => x"1e",
  4496 => x"c0",
  4497 => x"f6",
  4498 => x"ff",
  4499 => x"1e",
  4500 => x"d0",
  4501 => x"a6",
  4502 => x"1e",
  4503 => x"d0",
  4504 => x"66",
  4505 => x"1e",
  4506 => x"f8",
  4507 => x"e4",
  4508 => x"87",
  4509 => x"f0",
  4510 => x"8e",
  4511 => x"26",
  4512 => x"4f",
  4513 => x"1e",
  4514 => x"73",
  4515 => x"1e",
  4516 => x"72",
  4517 => x"9a",
  4518 => x"02",
  4519 => x"c0",
  4520 => x"e7",
  4521 => x"87",
  4522 => x"c0",
  4523 => x"48",
  4524 => x"c1",
  4525 => x"4b",
  4526 => x"72",
  4527 => x"a9",
  4528 => x"06",
  4529 => x"d1",
  4530 => x"87",
  4531 => x"72",
  4532 => x"82",
  4533 => x"06",
  4534 => x"c9",
  4535 => x"87",
  4536 => x"73",
  4537 => x"83",
  4538 => x"72",
  4539 => x"a9",
  4540 => x"01",
  4541 => x"f4",
  4542 => x"87",
  4543 => x"c3",
  4544 => x"87",
  4545 => x"c1",
  4546 => x"b2",
  4547 => x"3a",
  4548 => x"72",
  4549 => x"a9",
  4550 => x"03",
  4551 => x"89",
  4552 => x"73",
  4553 => x"80",
  4554 => x"07",
  4555 => x"c1",
  4556 => x"2a",
  4557 => x"2b",
  4558 => x"05",
  4559 => x"f3",
  4560 => x"87",
  4561 => x"26",
  4562 => x"4b",
  4563 => x"26",
  4564 => x"4f",
  4565 => x"1e",
  4566 => x"75",
  4567 => x"1e",
  4568 => x"c4",
  4569 => x"4d",
  4570 => x"71",
  4571 => x"b7",
  4572 => x"a1",
  4573 => x"04",
  4574 => x"ff",
  4575 => x"b9",
  4576 => x"c1",
  4577 => x"81",
  4578 => x"c3",
  4579 => x"bd",
  4580 => x"07",
  4581 => x"72",
  4582 => x"b7",
  4583 => x"a2",
  4584 => x"04",
  4585 => x"ff",
  4586 => x"ba",
  4587 => x"c1",
  4588 => x"82",
  4589 => x"c1",
  4590 => x"bd",
  4591 => x"07",
  4592 => x"fe",
  4593 => x"ee",
  4594 => x"87",
  4595 => x"c1",
  4596 => x"2d",
  4597 => x"04",
  4598 => x"ff",
  4599 => x"b8",
  4600 => x"c1",
  4601 => x"80",
  4602 => x"07",
  4603 => x"2d",
  4604 => x"04",
  4605 => x"ff",
  4606 => x"b9",
  4607 => x"c1",
  4608 => x"81",
  4609 => x"07",
  4610 => x"26",
  4611 => x"4d",
  4612 => x"26",
  4613 => x"4f",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;

