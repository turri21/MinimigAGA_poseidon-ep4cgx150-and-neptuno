library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"01",
     1 => x"da",
     2 => x"87",
     3 => x"04",
     4 => x"dd",
     5 => x"87",
     6 => x"0e",
     7 => x"58",
     8 => x"5e",
     9 => x"59",
    10 => x"5a",
    11 => x"0e",
    12 => x"27",
    13 => x"00",
    14 => x"00",
    15 => x"00",
    16 => x"2c",
    17 => x"0f",
    18 => x"26",
    19 => x"4a",
    20 => x"26",
    21 => x"49",
    22 => x"26",
    23 => x"48",
    24 => x"ff",
    25 => x"80",
    26 => x"26",
    27 => x"08",
    28 => x"4f",
    29 => x"27",
    30 => x"00",
    31 => x"00",
    32 => x"00",
    33 => x"2d",
    34 => x"4f",
    35 => x"27",
    36 => x"00",
    37 => x"00",
    38 => x"00",
    39 => x"29",
    40 => x"4f",
    41 => x"00",
    42 => x"fd",
    43 => x"87",
    44 => x"4f",
    45 => x"c1",
    46 => x"cc",
    47 => x"c8",
    48 => x"4e",
    49 => x"c9",
    50 => x"c0",
    51 => x"86",
    52 => x"c1",
    53 => x"cc",
    54 => x"c8",
    55 => x"49",
    56 => x"c1",
    57 => x"c2",
    58 => x"e4",
    59 => x"48",
    60 => x"89",
    61 => x"d0",
    62 => x"89",
    63 => x"03",
    64 => x"c0",
    65 => x"40",
    66 => x"40",
    67 => x"40",
    68 => x"40",
    69 => x"f6",
    70 => x"87",
    71 => x"d0",
    72 => x"81",
    73 => x"05",
    74 => x"c0",
    75 => x"50",
    76 => x"c1",
    77 => x"89",
    78 => x"05",
    79 => x"f9",
    80 => x"87",
    81 => x"c1",
    82 => x"c2",
    83 => x"e1",
    84 => x"4d",
    85 => x"c1",
    86 => x"c2",
    87 => x"e1",
    88 => x"4c",
    89 => x"74",
    90 => x"ad",
    91 => x"02",
    92 => x"c4",
    93 => x"87",
    94 => x"24",
    95 => x"0f",
    96 => x"f7",
    97 => x"87",
    98 => x"c1",
    99 => x"c0",
   100 => x"87",
   101 => x"c1",
   102 => x"c2",
   103 => x"e1",
   104 => x"4d",
   105 => x"c1",
   106 => x"c2",
   107 => x"e1",
   108 => x"4c",
   109 => x"74",
   110 => x"ad",
   111 => x"02",
   112 => x"c6",
   113 => x"87",
   114 => x"c4",
   115 => x"8c",
   116 => x"6c",
   117 => x"0f",
   118 => x"f5",
   119 => x"87",
   120 => x"00",
   121 => x"fd",
   122 => x"87",
   123 => x"1e",
   124 => x"73",
   125 => x"1e",
   126 => x"c2",
   127 => x"c0",
   128 => x"c0",
   129 => x"4b",
   130 => x"73",
   131 => x"0f",
   132 => x"c4",
   133 => x"87",
   134 => x"26",
   135 => x"4d",
   136 => x"26",
   137 => x"4c",
   138 => x"26",
   139 => x"4b",
   140 => x"26",
   141 => x"4f",
   142 => x"1e",
   143 => x"e5",
   144 => x"48",
   145 => x"c0",
   146 => x"e0",
   147 => x"50",
   148 => x"e5",
   149 => x"48",
   150 => x"c0",
   151 => x"e1",
   152 => x"50",
   153 => x"e5",
   154 => x"48",
   155 => x"c0",
   156 => x"e0",
   157 => x"50",
   158 => x"e5",
   159 => x"48",
   160 => x"c0",
   161 => x"e1",
   162 => x"50",
   163 => x"26",
   164 => x"4f",
   165 => x"1e",
   166 => x"73",
   167 => x"1e",
   168 => x"e5",
   169 => x"48",
   170 => x"c0",
   171 => x"e0",
   172 => x"50",
   173 => x"e5",
   174 => x"48",
   175 => x"c0",
   176 => x"e1",
   177 => x"50",
   178 => x"c5",
   179 => x"c4",
   180 => x"49",
   181 => x"c0",
   182 => x"f0",
   183 => x"e0",
   184 => x"87",
   185 => x"c0",
   186 => x"fc",
   187 => x"c0",
   188 => x"4b",
   189 => x"cf",
   190 => x"da",
   191 => x"87",
   192 => x"70",
   193 => x"98",
   194 => x"02",
   195 => x"c0",
   196 => x"f4",
   197 => x"87",
   198 => x"c0",
   199 => x"ff",
   200 => x"f0",
   201 => x"4b",
   202 => x"c4",
   203 => x"ed",
   204 => x"49",
   205 => x"c0",
   206 => x"f0",
   207 => x"c8",
   208 => x"87",
   209 => x"d5",
   210 => x"cd",
   211 => x"87",
   212 => x"70",
   213 => x"98",
   214 => x"02",
   215 => x"da",
   216 => x"87",
   217 => x"c3",
   218 => x"f0",
   219 => x"4b",
   220 => x"c2",
   221 => x"c0",
   222 => x"c0",
   223 => x"1e",
   224 => x"c4",
   225 => x"c5",
   226 => x"49",
   227 => x"c0",
   228 => x"ec",
   229 => x"ff",
   230 => x"87",
   231 => x"c4",
   232 => x"86",
   233 => x"70",
   234 => x"98",
   235 => x"02",
   236 => x"cc",
   237 => x"87",
   238 => x"fe",
   239 => x"ca",
   240 => x"87",
   241 => x"c7",
   242 => x"87",
   243 => x"c4",
   244 => x"d1",
   245 => x"49",
   246 => x"c0",
   247 => x"ef",
   248 => x"df",
   249 => x"87",
   250 => x"73",
   251 => x"49",
   252 => x"fe",
   253 => x"cf",
   254 => x"87",
   255 => x"fe",
   256 => x"f0",
   257 => x"87",
   258 => x"fe",
   259 => x"c5",
   260 => x"87",
   261 => x"38",
   262 => x"33",
   263 => x"32",
   264 => x"4f",
   265 => x"53",
   266 => x"44",
   267 => x"41",
   268 => x"42",
   269 => x"42",
   270 => x"49",
   271 => x"4e",
   272 => x"00",
   273 => x"55",
   274 => x"6e",
   275 => x"61",
   276 => x"62",
   277 => x"6c",
   278 => x"65",
   279 => x"20",
   280 => x"74",
   281 => x"6f",
   282 => x"20",
   283 => x"6c",
   284 => x"6f",
   285 => x"63",
   286 => x"61",
   287 => x"74",
   288 => x"65",
   289 => x"20",
   290 => x"70",
   291 => x"61",
   292 => x"72",
   293 => x"74",
   294 => x"69",
   295 => x"74",
   296 => x"69",
   297 => x"6f",
   298 => x"6e",
   299 => x"0a",
   300 => x"00",
   301 => x"48",
   302 => x"75",
   303 => x"6e",
   304 => x"74",
   305 => x"69",
   306 => x"6e",
   307 => x"67",
   308 => x"20",
   309 => x"66",
   310 => x"6f",
   311 => x"72",
   312 => x"20",
   313 => x"70",
   314 => x"61",
   315 => x"72",
   316 => x"74",
   317 => x"69",
   318 => x"74",
   319 => x"69",
   320 => x"6f",
   321 => x"6e",
   322 => x"0a",
   323 => x"00",
   324 => x"49",
   325 => x"6e",
   326 => x"69",
   327 => x"74",
   328 => x"69",
   329 => x"61",
   330 => x"6c",
   331 => x"69",
   332 => x"7a",
   333 => x"69",
   334 => x"6e",
   335 => x"67",
   336 => x"20",
   337 => x"53",
   338 => x"44",
   339 => x"20",
   340 => x"63",
   341 => x"61",
   342 => x"72",
   343 => x"64",
   344 => x"0a",
   345 => x"00",
   346 => x"1e",
   347 => x"e4",
   348 => x"86",
   349 => x"e1",
   350 => x"48",
   351 => x"c3",
   352 => x"ff",
   353 => x"50",
   354 => x"e1",
   355 => x"97",
   356 => x"bf",
   357 => x"48",
   358 => x"c4",
   359 => x"a6",
   360 => x"58",
   361 => x"6e",
   362 => x"49",
   363 => x"c3",
   364 => x"ff",
   365 => x"99",
   366 => x"e1",
   367 => x"48",
   368 => x"c3",
   369 => x"ff",
   370 => x"50",
   371 => x"c8",
   372 => x"31",
   373 => x"e1",
   374 => x"97",
   375 => x"bf",
   376 => x"48",
   377 => x"c8",
   378 => x"a6",
   379 => x"58",
   380 => x"c4",
   381 => x"66",
   382 => x"48",
   383 => x"c3",
   384 => x"ff",
   385 => x"98",
   386 => x"cc",
   387 => x"a6",
   388 => x"58",
   389 => x"c8",
   390 => x"66",
   391 => x"b1",
   392 => x"e1",
   393 => x"48",
   394 => x"c3",
   395 => x"ff",
   396 => x"50",
   397 => x"c8",
   398 => x"31",
   399 => x"e1",
   400 => x"97",
   401 => x"bf",
   402 => x"48",
   403 => x"d0",
   404 => x"a6",
   405 => x"58",
   406 => x"cc",
   407 => x"66",
   408 => x"48",
   409 => x"c3",
   410 => x"ff",
   411 => x"98",
   412 => x"d4",
   413 => x"a6",
   414 => x"58",
   415 => x"d0",
   416 => x"66",
   417 => x"b1",
   418 => x"e1",
   419 => x"48",
   420 => x"c3",
   421 => x"ff",
   422 => x"50",
   423 => x"c8",
   424 => x"31",
   425 => x"e1",
   426 => x"97",
   427 => x"bf",
   428 => x"48",
   429 => x"d8",
   430 => x"a6",
   431 => x"58",
   432 => x"d4",
   433 => x"66",
   434 => x"48",
   435 => x"c3",
   436 => x"ff",
   437 => x"98",
   438 => x"dc",
   439 => x"a6",
   440 => x"58",
   441 => x"d8",
   442 => x"66",
   443 => x"b1",
   444 => x"71",
   445 => x"48",
   446 => x"e4",
   447 => x"8e",
   448 => x"26",
   449 => x"4f",
   450 => x"0e",
   451 => x"5e",
   452 => x"5b",
   453 => x"5c",
   454 => x"0e",
   455 => x"1e",
   456 => x"71",
   457 => x"4a",
   458 => x"72",
   459 => x"49",
   460 => x"c3",
   461 => x"ff",
   462 => x"99",
   463 => x"e1",
   464 => x"09",
   465 => x"97",
   466 => x"79",
   467 => x"09",
   468 => x"c1",
   469 => x"c2",
   470 => x"e4",
   471 => x"bf",
   472 => x"05",
   473 => x"c8",
   474 => x"87",
   475 => x"d0",
   476 => x"66",
   477 => x"48",
   478 => x"c9",
   479 => x"30",
   480 => x"d4",
   481 => x"a6",
   482 => x"58",
   483 => x"d0",
   484 => x"66",
   485 => x"49",
   486 => x"d8",
   487 => x"29",
   488 => x"c3",
   489 => x"ff",
   490 => x"99",
   491 => x"e1",
   492 => x"09",
   493 => x"97",
   494 => x"79",
   495 => x"09",
   496 => x"d0",
   497 => x"66",
   498 => x"49",
   499 => x"d0",
   500 => x"29",
   501 => x"c3",
   502 => x"ff",
   503 => x"99",
   504 => x"e1",
   505 => x"09",
   506 => x"97",
   507 => x"79",
   508 => x"09",
   509 => x"d0",
   510 => x"66",
   511 => x"49",
   512 => x"c8",
   513 => x"29",
   514 => x"c3",
   515 => x"ff",
   516 => x"99",
   517 => x"e1",
   518 => x"09",
   519 => x"97",
   520 => x"79",
   521 => x"09",
   522 => x"d0",
   523 => x"66",
   524 => x"49",
   525 => x"c3",
   526 => x"ff",
   527 => x"99",
   528 => x"e1",
   529 => x"09",
   530 => x"97",
   531 => x"79",
   532 => x"09",
   533 => x"72",
   534 => x"49",
   535 => x"d0",
   536 => x"29",
   537 => x"c3",
   538 => x"ff",
   539 => x"99",
   540 => x"e1",
   541 => x"09",
   542 => x"97",
   543 => x"79",
   544 => x"09",
   545 => x"97",
   546 => x"bf",
   547 => x"48",
   548 => x"c4",
   549 => x"a6",
   550 => x"58",
   551 => x"6e",
   552 => x"4b",
   553 => x"c3",
   554 => x"ff",
   555 => x"9b",
   556 => x"c9",
   557 => x"f0",
   558 => x"ff",
   559 => x"4c",
   560 => x"c3",
   561 => x"ff",
   562 => x"ab",
   563 => x"05",
   564 => x"dc",
   565 => x"87",
   566 => x"e1",
   567 => x"48",
   568 => x"c3",
   569 => x"ff",
   570 => x"50",
   571 => x"e1",
   572 => x"97",
   573 => x"bf",
   574 => x"48",
   575 => x"c4",
   576 => x"a6",
   577 => x"58",
   578 => x"6e",
   579 => x"4b",
   580 => x"c3",
   581 => x"ff",
   582 => x"9b",
   583 => x"c1",
   584 => x"8c",
   585 => x"02",
   586 => x"c6",
   587 => x"87",
   588 => x"c3",
   589 => x"ff",
   590 => x"ab",
   591 => x"02",
   592 => x"e4",
   593 => x"87",
   594 => x"73",
   595 => x"4a",
   596 => x"c4",
   597 => x"b7",
   598 => x"2a",
   599 => x"c0",
   600 => x"f0",
   601 => x"a2",
   602 => x"49",
   603 => x"c0",
   604 => x"e9",
   605 => x"f0",
   606 => x"87",
   607 => x"73",
   608 => x"4a",
   609 => x"cf",
   610 => x"9a",
   611 => x"c0",
   612 => x"f0",
   613 => x"a2",
   614 => x"49",
   615 => x"c0",
   616 => x"e9",
   617 => x"e4",
   618 => x"87",
   619 => x"73",
   620 => x"48",
   621 => x"26",
   622 => x"c2",
   623 => x"87",
   624 => x"26",
   625 => x"4d",
   626 => x"26",
   627 => x"4c",
   628 => x"26",
   629 => x"4b",
   630 => x"26",
   631 => x"4f",
   632 => x"1e",
   633 => x"c0",
   634 => x"49",
   635 => x"e1",
   636 => x"48",
   637 => x"c3",
   638 => x"ff",
   639 => x"50",
   640 => x"c1",
   641 => x"81",
   642 => x"c3",
   643 => x"c8",
   644 => x"b7",
   645 => x"a9",
   646 => x"04",
   647 => x"f2",
   648 => x"87",
   649 => x"26",
   650 => x"4f",
   651 => x"1e",
   652 => x"73",
   653 => x"1e",
   654 => x"e8",
   655 => x"87",
   656 => x"c4",
   657 => x"f8",
   658 => x"df",
   659 => x"4b",
   660 => x"c0",
   661 => x"1e",
   662 => x"c0",
   663 => x"ff",
   664 => x"f0",
   665 => x"c1",
   666 => x"f7",
   667 => x"49",
   668 => x"fc",
   669 => x"e3",
   670 => x"87",
   671 => x"c4",
   672 => x"86",
   673 => x"c1",
   674 => x"a8",
   675 => x"05",
   676 => x"c0",
   677 => x"e8",
   678 => x"87",
   679 => x"e1",
   680 => x"48",
   681 => x"c3",
   682 => x"ff",
   683 => x"50",
   684 => x"c1",
   685 => x"c0",
   686 => x"c0",
   687 => x"c0",
   688 => x"c0",
   689 => x"c0",
   690 => x"1e",
   691 => x"c0",
   692 => x"e1",
   693 => x"f0",
   694 => x"c1",
   695 => x"e9",
   696 => x"49",
   697 => x"fc",
   698 => x"c6",
   699 => x"87",
   700 => x"c4",
   701 => x"86",
   702 => x"70",
   703 => x"98",
   704 => x"05",
   705 => x"c9",
   706 => x"87",
   707 => x"e1",
   708 => x"48",
   709 => x"c3",
   710 => x"ff",
   711 => x"50",
   712 => x"c1",
   713 => x"48",
   714 => x"cb",
   715 => x"87",
   716 => x"fe",
   717 => x"e9",
   718 => x"87",
   719 => x"c1",
   720 => x"8b",
   721 => x"05",
   722 => x"fe",
   723 => x"ff",
   724 => x"87",
   725 => x"c0",
   726 => x"48",
   727 => x"fe",
   728 => x"da",
   729 => x"87",
   730 => x"43",
   731 => x"4d",
   732 => x"44",
   733 => x"34",
   734 => x"31",
   735 => x"20",
   736 => x"25",
   737 => x"64",
   738 => x"0a",
   739 => x"00",
   740 => x"43",
   741 => x"4d",
   742 => x"44",
   743 => x"35",
   744 => x"35",
   745 => x"20",
   746 => x"25",
   747 => x"64",
   748 => x"0a",
   749 => x"00",
   750 => x"43",
   751 => x"4d",
   752 => x"44",
   753 => x"34",
   754 => x"31",
   755 => x"20",
   756 => x"25",
   757 => x"64",
   758 => x"0a",
   759 => x"00",
   760 => x"43",
   761 => x"4d",
   762 => x"44",
   763 => x"35",
   764 => x"35",
   765 => x"20",
   766 => x"25",
   767 => x"64",
   768 => x"0a",
   769 => x"00",
   770 => x"69",
   771 => x"6e",
   772 => x"69",
   773 => x"74",
   774 => x"20",
   775 => x"25",
   776 => x"64",
   777 => x"0a",
   778 => x"20",
   779 => x"20",
   780 => x"00",
   781 => x"69",
   782 => x"6e",
   783 => x"69",
   784 => x"74",
   785 => x"20",
   786 => x"25",
   787 => x"64",
   788 => x"0a",
   789 => x"20",
   790 => x"20",
   791 => x"00",
   792 => x"43",
   793 => x"6d",
   794 => x"64",
   795 => x"5f",
   796 => x"69",
   797 => x"6e",
   798 => x"69",
   799 => x"74",
   800 => x"0a",
   801 => x"00",
   802 => x"43",
   803 => x"4d",
   804 => x"44",
   805 => x"38",
   806 => x"5f",
   807 => x"34",
   808 => x"20",
   809 => x"72",
   810 => x"65",
   811 => x"73",
   812 => x"70",
   813 => x"6f",
   814 => x"6e",
   815 => x"73",
   816 => x"65",
   817 => x"3a",
   818 => x"20",
   819 => x"25",
   820 => x"64",
   821 => x"0a",
   822 => x"00",
   823 => x"43",
   824 => x"4d",
   825 => x"44",
   826 => x"35",
   827 => x"38",
   828 => x"20",
   829 => x"25",
   830 => x"64",
   831 => x"0a",
   832 => x"20",
   833 => x"20",
   834 => x"00",
   835 => x"43",
   836 => x"4d",
   837 => x"44",
   838 => x"35",
   839 => x"38",
   840 => x"5f",
   841 => x"32",
   842 => x"20",
   843 => x"25",
   844 => x"64",
   845 => x"0a",
   846 => x"20",
   847 => x"20",
   848 => x"00",
   849 => x"43",
   850 => x"4d",
   851 => x"44",
   852 => x"35",
   853 => x"38",
   854 => x"20",
   855 => x"25",
   856 => x"64",
   857 => x"0a",
   858 => x"20",
   859 => x"20",
   860 => x"00",
   861 => x"53",
   862 => x"44",
   863 => x"48",
   864 => x"43",
   865 => x"20",
   866 => x"49",
   867 => x"6e",
   868 => x"69",
   869 => x"74",
   870 => x"69",
   871 => x"61",
   872 => x"6c",
   873 => x"69",
   874 => x"7a",
   875 => x"61",
   876 => x"74",
   877 => x"69",
   878 => x"6f",
   879 => x"6e",
   880 => x"20",
   881 => x"65",
   882 => x"72",
   883 => x"72",
   884 => x"6f",
   885 => x"72",
   886 => x"21",
   887 => x"0a",
   888 => x"00",
   889 => x"63",
   890 => x"6d",
   891 => x"64",
   892 => x"5f",
   893 => x"43",
   894 => x"4d",
   895 => x"44",
   896 => x"38",
   897 => x"20",
   898 => x"72",
   899 => x"65",
   900 => x"73",
   901 => x"70",
   902 => x"6f",
   903 => x"6e",
   904 => x"73",
   905 => x"65",
   906 => x"3a",
   907 => x"20",
   908 => x"25",
   909 => x"64",
   910 => x"0a",
   911 => x"00",
   912 => x"52",
   913 => x"65",
   914 => x"61",
   915 => x"64",
   916 => x"20",
   917 => x"63",
   918 => x"6f",
   919 => x"6d",
   920 => x"6d",
   921 => x"61",
   922 => x"6e",
   923 => x"64",
   924 => x"20",
   925 => x"66",
   926 => x"61",
   927 => x"69",
   928 => x"6c",
   929 => x"65",
   930 => x"64",
   931 => x"20",
   932 => x"61",
   933 => x"74",
   934 => x"20",
   935 => x"25",
   936 => x"64",
   937 => x"20",
   938 => x"28",
   939 => x"25",
   940 => x"64",
   941 => x"29",
   942 => x"0a",
   943 => x"00",
   944 => x"1e",
   945 => x"73",
   946 => x"1e",
   947 => x"e1",
   948 => x"48",
   949 => x"c3",
   950 => x"ff",
   951 => x"50",
   952 => x"cc",
   953 => x"d8",
   954 => x"49",
   955 => x"c0",
   956 => x"e4",
   957 => x"da",
   958 => x"87",
   959 => x"d3",
   960 => x"4b",
   961 => x"c0",
   962 => x"1e",
   963 => x"c0",
   964 => x"ff",
   965 => x"f0",
   966 => x"c1",
   967 => x"c1",
   968 => x"49",
   969 => x"f7",
   970 => x"f6",
   971 => x"87",
   972 => x"c4",
   973 => x"86",
   974 => x"70",
   975 => x"98",
   976 => x"05",
   977 => x"c9",
   978 => x"87",
   979 => x"e1",
   980 => x"48",
   981 => x"c3",
   982 => x"ff",
   983 => x"50",
   984 => x"c1",
   985 => x"48",
   986 => x"cb",
   987 => x"87",
   988 => x"fa",
   989 => x"d9",
   990 => x"87",
   991 => x"c1",
   992 => x"8b",
   993 => x"05",
   994 => x"ff",
   995 => x"dc",
   996 => x"87",
   997 => x"c0",
   998 => x"48",
   999 => x"fa",
  1000 => x"ca",
  1001 => x"87",
  1002 => x"1e",
  1003 => x"73",
  1004 => x"1e",
  1005 => x"1e",
  1006 => x"fa",
  1007 => x"c7",
  1008 => x"87",
  1009 => x"c6",
  1010 => x"ea",
  1011 => x"1e",
  1012 => x"c0",
  1013 => x"e1",
  1014 => x"f0",
  1015 => x"c1",
  1016 => x"c8",
  1017 => x"49",
  1018 => x"f7",
  1019 => x"c5",
  1020 => x"87",
  1021 => x"70",
  1022 => x"4b",
  1023 => x"73",
  1024 => x"1e",
  1025 => x"cd",
  1026 => x"f9",
  1027 => x"49",
  1028 => x"c0",
  1029 => x"f0",
  1030 => x"e0",
  1031 => x"87",
  1032 => x"c8",
  1033 => x"86",
  1034 => x"c1",
  1035 => x"ab",
  1036 => x"02",
  1037 => x"c8",
  1038 => x"87",
  1039 => x"fe",
  1040 => x"de",
  1041 => x"87",
  1042 => x"c0",
  1043 => x"48",
  1044 => x"c1",
  1045 => x"ff",
  1046 => x"87",
  1047 => x"f5",
  1048 => x"c0",
  1049 => x"87",
  1050 => x"70",
  1051 => x"49",
  1052 => x"cf",
  1053 => x"ff",
  1054 => x"ff",
  1055 => x"99",
  1056 => x"c6",
  1057 => x"ea",
  1058 => x"a9",
  1059 => x"02",
  1060 => x"c8",
  1061 => x"87",
  1062 => x"fe",
  1063 => x"c7",
  1064 => x"87",
  1065 => x"c0",
  1066 => x"48",
  1067 => x"c1",
  1068 => x"e8",
  1069 => x"87",
  1070 => x"e1",
  1071 => x"48",
  1072 => x"c3",
  1073 => x"ff",
  1074 => x"50",
  1075 => x"c0",
  1076 => x"f1",
  1077 => x"4b",
  1078 => x"f9",
  1079 => x"d2",
  1080 => x"87",
  1081 => x"70",
  1082 => x"98",
  1083 => x"02",
  1084 => x"c1",
  1085 => x"c6",
  1086 => x"87",
  1087 => x"c0",
  1088 => x"1e",
  1089 => x"c0",
  1090 => x"ff",
  1091 => x"f0",
  1092 => x"c1",
  1093 => x"fa",
  1094 => x"49",
  1095 => x"f5",
  1096 => x"f8",
  1097 => x"87",
  1098 => x"c4",
  1099 => x"86",
  1100 => x"70",
  1101 => x"98",
  1102 => x"05",
  1103 => x"c0",
  1104 => x"f3",
  1105 => x"87",
  1106 => x"e1",
  1107 => x"48",
  1108 => x"c3",
  1109 => x"ff",
  1110 => x"50",
  1111 => x"e1",
  1112 => x"97",
  1113 => x"bf",
  1114 => x"48",
  1115 => x"c4",
  1116 => x"a6",
  1117 => x"58",
  1118 => x"6e",
  1119 => x"49",
  1120 => x"c3",
  1121 => x"ff",
  1122 => x"99",
  1123 => x"e1",
  1124 => x"48",
  1125 => x"c3",
  1126 => x"ff",
  1127 => x"50",
  1128 => x"e1",
  1129 => x"48",
  1130 => x"c3",
  1131 => x"ff",
  1132 => x"50",
  1133 => x"e1",
  1134 => x"48",
  1135 => x"c3",
  1136 => x"ff",
  1137 => x"50",
  1138 => x"e1",
  1139 => x"48",
  1140 => x"c3",
  1141 => x"ff",
  1142 => x"50",
  1143 => x"c1",
  1144 => x"c0",
  1145 => x"99",
  1146 => x"02",
  1147 => x"c4",
  1148 => x"87",
  1149 => x"c1",
  1150 => x"48",
  1151 => x"d5",
  1152 => x"87",
  1153 => x"c0",
  1154 => x"48",
  1155 => x"d1",
  1156 => x"87",
  1157 => x"c2",
  1158 => x"ab",
  1159 => x"05",
  1160 => x"c4",
  1161 => x"87",
  1162 => x"c0",
  1163 => x"48",
  1164 => x"c8",
  1165 => x"87",
  1166 => x"c1",
  1167 => x"8b",
  1168 => x"05",
  1169 => x"fe",
  1170 => x"e2",
  1171 => x"87",
  1172 => x"c0",
  1173 => x"48",
  1174 => x"26",
  1175 => x"f7",
  1176 => x"da",
  1177 => x"87",
  1178 => x"1e",
  1179 => x"73",
  1180 => x"1e",
  1181 => x"c1",
  1182 => x"c2",
  1183 => x"e4",
  1184 => x"48",
  1185 => x"c1",
  1186 => x"78",
  1187 => x"e9",
  1188 => x"48",
  1189 => x"c3",
  1190 => x"ef",
  1191 => x"50",
  1192 => x"c7",
  1193 => x"4b",
  1194 => x"e5",
  1195 => x"48",
  1196 => x"c3",
  1197 => x"50",
  1198 => x"f7",
  1199 => x"c7",
  1200 => x"87",
  1201 => x"e5",
  1202 => x"48",
  1203 => x"c2",
  1204 => x"50",
  1205 => x"e1",
  1206 => x"48",
  1207 => x"c3",
  1208 => x"ff",
  1209 => x"50",
  1210 => x"c0",
  1211 => x"1e",
  1212 => x"c0",
  1213 => x"e5",
  1214 => x"d0",
  1215 => x"c1",
  1216 => x"c0",
  1217 => x"49",
  1218 => x"f3",
  1219 => x"fd",
  1220 => x"87",
  1221 => x"c4",
  1222 => x"86",
  1223 => x"c1",
  1224 => x"a8",
  1225 => x"05",
  1226 => x"c2",
  1227 => x"87",
  1228 => x"c1",
  1229 => x"4b",
  1230 => x"c2",
  1231 => x"ab",
  1232 => x"05",
  1233 => x"c5",
  1234 => x"87",
  1235 => x"c0",
  1236 => x"48",
  1237 => x"c0",
  1238 => x"f1",
  1239 => x"87",
  1240 => x"c1",
  1241 => x"8b",
  1242 => x"05",
  1243 => x"ff",
  1244 => x"cc",
  1245 => x"87",
  1246 => x"fc",
  1247 => x"c9",
  1248 => x"87",
  1249 => x"c1",
  1250 => x"c2",
  1251 => x"e8",
  1252 => x"58",
  1253 => x"c1",
  1254 => x"c2",
  1255 => x"e4",
  1256 => x"bf",
  1257 => x"05",
  1258 => x"cd",
  1259 => x"87",
  1260 => x"c1",
  1261 => x"1e",
  1262 => x"c0",
  1263 => x"ff",
  1264 => x"f0",
  1265 => x"c1",
  1266 => x"d0",
  1267 => x"49",
  1268 => x"f3",
  1269 => x"cb",
  1270 => x"87",
  1271 => x"c4",
  1272 => x"86",
  1273 => x"e1",
  1274 => x"48",
  1275 => x"c3",
  1276 => x"ff",
  1277 => x"50",
  1278 => x"e5",
  1279 => x"48",
  1280 => x"c3",
  1281 => x"50",
  1282 => x"e1",
  1283 => x"48",
  1284 => x"c3",
  1285 => x"ff",
  1286 => x"50",
  1287 => x"c1",
  1288 => x"48",
  1289 => x"f5",
  1290 => x"e8",
  1291 => x"87",
  1292 => x"0e",
  1293 => x"5e",
  1294 => x"5b",
  1295 => x"5c",
  1296 => x"5d",
  1297 => x"0e",
  1298 => x"1e",
  1299 => x"71",
  1300 => x"4a",
  1301 => x"c0",
  1302 => x"4d",
  1303 => x"e1",
  1304 => x"48",
  1305 => x"c3",
  1306 => x"ff",
  1307 => x"50",
  1308 => x"e5",
  1309 => x"48",
  1310 => x"c2",
  1311 => x"50",
  1312 => x"e9",
  1313 => x"48",
  1314 => x"c7",
  1315 => x"50",
  1316 => x"e1",
  1317 => x"48",
  1318 => x"c3",
  1319 => x"ff",
  1320 => x"50",
  1321 => x"72",
  1322 => x"1e",
  1323 => x"c0",
  1324 => x"ff",
  1325 => x"f0",
  1326 => x"c1",
  1327 => x"d1",
  1328 => x"49",
  1329 => x"f2",
  1330 => x"ce",
  1331 => x"87",
  1332 => x"c4",
  1333 => x"86",
  1334 => x"70",
  1335 => x"98",
  1336 => x"05",
  1337 => x"c1",
  1338 => x"c9",
  1339 => x"87",
  1340 => x"c5",
  1341 => x"ee",
  1342 => x"cd",
  1343 => x"df",
  1344 => x"4b",
  1345 => x"e1",
  1346 => x"48",
  1347 => x"c3",
  1348 => x"ff",
  1349 => x"50",
  1350 => x"e1",
  1351 => x"97",
  1352 => x"bf",
  1353 => x"48",
  1354 => x"c4",
  1355 => x"a6",
  1356 => x"58",
  1357 => x"6e",
  1358 => x"49",
  1359 => x"c3",
  1360 => x"ff",
  1361 => x"99",
  1362 => x"c3",
  1363 => x"fe",
  1364 => x"a9",
  1365 => x"05",
  1366 => x"de",
  1367 => x"87",
  1368 => x"c0",
  1369 => x"4c",
  1370 => x"ef",
  1371 => x"fd",
  1372 => x"87",
  1373 => x"d4",
  1374 => x"66",
  1375 => x"08",
  1376 => x"78",
  1377 => x"08",
  1378 => x"d4",
  1379 => x"66",
  1380 => x"48",
  1381 => x"c4",
  1382 => x"80",
  1383 => x"d8",
  1384 => x"a6",
  1385 => x"58",
  1386 => x"c1",
  1387 => x"84",
  1388 => x"c2",
  1389 => x"c0",
  1390 => x"b7",
  1391 => x"ac",
  1392 => x"04",
  1393 => x"e7",
  1394 => x"87",
  1395 => x"c1",
  1396 => x"4b",
  1397 => x"4d",
  1398 => x"c1",
  1399 => x"8b",
  1400 => x"05",
  1401 => x"ff",
  1402 => x"c5",
  1403 => x"87",
  1404 => x"e1",
  1405 => x"48",
  1406 => x"c3",
  1407 => x"ff",
  1408 => x"50",
  1409 => x"e5",
  1410 => x"48",
  1411 => x"c3",
  1412 => x"50",
  1413 => x"75",
  1414 => x"48",
  1415 => x"26",
  1416 => x"f3",
  1417 => x"e5",
  1418 => x"87",
  1419 => x"1e",
  1420 => x"73",
  1421 => x"1e",
  1422 => x"71",
  1423 => x"4b",
  1424 => x"73",
  1425 => x"49",
  1426 => x"d8",
  1427 => x"29",
  1428 => x"c3",
  1429 => x"ff",
  1430 => x"99",
  1431 => x"73",
  1432 => x"4a",
  1433 => x"c8",
  1434 => x"2a",
  1435 => x"cf",
  1436 => x"fc",
  1437 => x"c0",
  1438 => x"9a",
  1439 => x"72",
  1440 => x"b1",
  1441 => x"73",
  1442 => x"4a",
  1443 => x"c8",
  1444 => x"32",
  1445 => x"c0",
  1446 => x"ff",
  1447 => x"f0",
  1448 => x"c0",
  1449 => x"c0",
  1450 => x"9a",
  1451 => x"72",
  1452 => x"b1",
  1453 => x"73",
  1454 => x"4a",
  1455 => x"d8",
  1456 => x"32",
  1457 => x"ff",
  1458 => x"c0",
  1459 => x"c0",
  1460 => x"c0",
  1461 => x"c0",
  1462 => x"9a",
  1463 => x"72",
  1464 => x"b1",
  1465 => x"71",
  1466 => x"48",
  1467 => x"c4",
  1468 => x"87",
  1469 => x"26",
  1470 => x"4d",
  1471 => x"26",
  1472 => x"4c",
  1473 => x"26",
  1474 => x"4b",
  1475 => x"26",
  1476 => x"4f",
  1477 => x"1e",
  1478 => x"73",
  1479 => x"1e",
  1480 => x"71",
  1481 => x"4b",
  1482 => x"73",
  1483 => x"49",
  1484 => x"c8",
  1485 => x"29",
  1486 => x"c3",
  1487 => x"ff",
  1488 => x"99",
  1489 => x"73",
  1490 => x"4a",
  1491 => x"c8",
  1492 => x"32",
  1493 => x"cf",
  1494 => x"fc",
  1495 => x"c0",
  1496 => x"9a",
  1497 => x"72",
  1498 => x"b1",
  1499 => x"71",
  1500 => x"48",
  1501 => x"e2",
  1502 => x"87",
  1503 => x"0e",
  1504 => x"5e",
  1505 => x"5b",
  1506 => x"5c",
  1507 => x"0e",
  1508 => x"71",
  1509 => x"4b",
  1510 => x"c0",
  1511 => x"4c",
  1512 => x"d0",
  1513 => x"66",
  1514 => x"48",
  1515 => x"c0",
  1516 => x"b7",
  1517 => x"a8",
  1518 => x"06",
  1519 => x"c0",
  1520 => x"e3",
  1521 => x"87",
  1522 => x"13",
  1523 => x"4a",
  1524 => x"cc",
  1525 => x"66",
  1526 => x"97",
  1527 => x"bf",
  1528 => x"49",
  1529 => x"cc",
  1530 => x"66",
  1531 => x"48",
  1532 => x"c1",
  1533 => x"80",
  1534 => x"d0",
  1535 => x"a6",
  1536 => x"58",
  1537 => x"71",
  1538 => x"b7",
  1539 => x"aa",
  1540 => x"02",
  1541 => x"c4",
  1542 => x"87",
  1543 => x"c1",
  1544 => x"48",
  1545 => x"cc",
  1546 => x"87",
  1547 => x"c1",
  1548 => x"84",
  1549 => x"d0",
  1550 => x"66",
  1551 => x"b7",
  1552 => x"ac",
  1553 => x"04",
  1554 => x"ff",
  1555 => x"dd",
  1556 => x"87",
  1557 => x"c0",
  1558 => x"48",
  1559 => x"c2",
  1560 => x"87",
  1561 => x"26",
  1562 => x"4d",
  1563 => x"26",
  1564 => x"4c",
  1565 => x"26",
  1566 => x"4b",
  1567 => x"26",
  1568 => x"4f",
  1569 => x"0e",
  1570 => x"5e",
  1571 => x"5b",
  1572 => x"5c",
  1573 => x"5d",
  1574 => x"0e",
  1575 => x"c1",
  1576 => x"cb",
  1577 => x"e6",
  1578 => x"48",
  1579 => x"ff",
  1580 => x"78",
  1581 => x"c1",
  1582 => x"ca",
  1583 => x"f6",
  1584 => x"48",
  1585 => x"c0",
  1586 => x"78",
  1587 => x"c0",
  1588 => x"e6",
  1589 => x"d6",
  1590 => x"49",
  1591 => x"da",
  1592 => x"df",
  1593 => x"87",
  1594 => x"c1",
  1595 => x"c2",
  1596 => x"ee",
  1597 => x"1e",
  1598 => x"c0",
  1599 => x"49",
  1600 => x"fb",
  1601 => x"c9",
  1602 => x"87",
  1603 => x"c4",
  1604 => x"86",
  1605 => x"70",
  1606 => x"98",
  1607 => x"05",
  1608 => x"c5",
  1609 => x"87",
  1610 => x"c0",
  1611 => x"48",
  1612 => x"cb",
  1613 => x"c1",
  1614 => x"87",
  1615 => x"c0",
  1616 => x"4b",
  1617 => x"c1",
  1618 => x"cb",
  1619 => x"e2",
  1620 => x"48",
  1621 => x"c1",
  1622 => x"78",
  1623 => x"c8",
  1624 => x"1e",
  1625 => x"c0",
  1626 => x"e6",
  1627 => x"e3",
  1628 => x"1e",
  1629 => x"c1",
  1630 => x"c3",
  1631 => x"e4",
  1632 => x"49",
  1633 => x"fd",
  1634 => x"fb",
  1635 => x"87",
  1636 => x"c8",
  1637 => x"86",
  1638 => x"70",
  1639 => x"98",
  1640 => x"05",
  1641 => x"c6",
  1642 => x"87",
  1643 => x"c1",
  1644 => x"cb",
  1645 => x"e2",
  1646 => x"48",
  1647 => x"c0",
  1648 => x"78",
  1649 => x"c8",
  1650 => x"1e",
  1651 => x"c0",
  1652 => x"e6",
  1653 => x"ec",
  1654 => x"1e",
  1655 => x"c1",
  1656 => x"c4",
  1657 => x"c0",
  1658 => x"49",
  1659 => x"fd",
  1660 => x"e1",
  1661 => x"87",
  1662 => x"c8",
  1663 => x"86",
  1664 => x"70",
  1665 => x"98",
  1666 => x"05",
  1667 => x"c6",
  1668 => x"87",
  1669 => x"c1",
  1670 => x"cb",
  1671 => x"e2",
  1672 => x"48",
  1673 => x"c0",
  1674 => x"78",
  1675 => x"c8",
  1676 => x"1e",
  1677 => x"c0",
  1678 => x"e6",
  1679 => x"f5",
  1680 => x"1e",
  1681 => x"c1",
  1682 => x"c4",
  1683 => x"c0",
  1684 => x"49",
  1685 => x"fd",
  1686 => x"c7",
  1687 => x"87",
  1688 => x"c8",
  1689 => x"86",
  1690 => x"70",
  1691 => x"98",
  1692 => x"05",
  1693 => x"c5",
  1694 => x"87",
  1695 => x"c0",
  1696 => x"48",
  1697 => x"c9",
  1698 => x"ec",
  1699 => x"87",
  1700 => x"c1",
  1701 => x"cb",
  1702 => x"e2",
  1703 => x"bf",
  1704 => x"1e",
  1705 => x"c0",
  1706 => x"e6",
  1707 => x"fe",
  1708 => x"1e",
  1709 => x"c0",
  1710 => x"e5",
  1711 => x"f7",
  1712 => x"87",
  1713 => x"c8",
  1714 => x"86",
  1715 => x"c1",
  1716 => x"cb",
  1717 => x"e2",
  1718 => x"bf",
  1719 => x"02",
  1720 => x"c1",
  1721 => x"f4",
  1722 => x"87",
  1723 => x"c1",
  1724 => x"c2",
  1725 => x"ee",
  1726 => x"4d",
  1727 => x"48",
  1728 => x"c6",
  1729 => x"fe",
  1730 => x"a0",
  1731 => x"4c",
  1732 => x"c8",
  1733 => x"c0",
  1734 => x"1e",
  1735 => x"70",
  1736 => x"49",
  1737 => x"d8",
  1738 => x"f6",
  1739 => x"87",
  1740 => x"c4",
  1741 => x"86",
  1742 => x"c8",
  1743 => x"a4",
  1744 => x"49",
  1745 => x"69",
  1746 => x"4b",
  1747 => x"c1",
  1748 => x"ca",
  1749 => x"ec",
  1750 => x"9f",
  1751 => x"bf",
  1752 => x"49",
  1753 => x"c5",
  1754 => x"d6",
  1755 => x"ea",
  1756 => x"a9",
  1757 => x"05",
  1758 => x"c0",
  1759 => x"cc",
  1760 => x"87",
  1761 => x"c8",
  1762 => x"a4",
  1763 => x"4a",
  1764 => x"6a",
  1765 => x"49",
  1766 => x"fa",
  1767 => x"e2",
  1768 => x"87",
  1769 => x"70",
  1770 => x"4b",
  1771 => x"db",
  1772 => x"87",
  1773 => x"c7",
  1774 => x"fe",
  1775 => x"a5",
  1776 => x"49",
  1777 => x"9f",
  1778 => x"69",
  1779 => x"49",
  1780 => x"ca",
  1781 => x"e9",
  1782 => x"d5",
  1783 => x"a9",
  1784 => x"02",
  1785 => x"c0",
  1786 => x"cc",
  1787 => x"87",
  1788 => x"c0",
  1789 => x"e4",
  1790 => x"d3",
  1791 => x"49",
  1792 => x"d7",
  1793 => x"d6",
  1794 => x"87",
  1795 => x"c0",
  1796 => x"48",
  1797 => x"c8",
  1798 => x"c8",
  1799 => x"87",
  1800 => x"73",
  1801 => x"1e",
  1802 => x"c0",
  1803 => x"e4",
  1804 => x"f1",
  1805 => x"1e",
  1806 => x"c0",
  1807 => x"e4",
  1808 => x"d6",
  1809 => x"87",
  1810 => x"c1",
  1811 => x"c2",
  1812 => x"ee",
  1813 => x"1e",
  1814 => x"73",
  1815 => x"49",
  1816 => x"f7",
  1817 => x"f1",
  1818 => x"87",
  1819 => x"cc",
  1820 => x"86",
  1821 => x"70",
  1822 => x"98",
  1823 => x"05",
  1824 => x"c0",
  1825 => x"c5",
  1826 => x"87",
  1827 => x"c0",
  1828 => x"48",
  1829 => x"c7",
  1830 => x"e8",
  1831 => x"87",
  1832 => x"c0",
  1833 => x"e5",
  1834 => x"c9",
  1835 => x"49",
  1836 => x"d6",
  1837 => x"ea",
  1838 => x"87",
  1839 => x"c8",
  1840 => x"c0",
  1841 => x"1e",
  1842 => x"c1",
  1843 => x"c2",
  1844 => x"ee",
  1845 => x"49",
  1846 => x"d7",
  1847 => x"c9",
  1848 => x"87",
  1849 => x"c0",
  1850 => x"e7",
  1851 => x"d1",
  1852 => x"1e",
  1853 => x"c0",
  1854 => x"e3",
  1855 => x"e7",
  1856 => x"87",
  1857 => x"c8",
  1858 => x"1e",
  1859 => x"c0",
  1860 => x"e7",
  1861 => x"e9",
  1862 => x"1e",
  1863 => x"c1",
  1864 => x"c4",
  1865 => x"c0",
  1866 => x"49",
  1867 => x"fa",
  1868 => x"d1",
  1869 => x"87",
  1870 => x"d0",
  1871 => x"86",
  1872 => x"70",
  1873 => x"98",
  1874 => x"05",
  1875 => x"c0",
  1876 => x"c9",
  1877 => x"87",
  1878 => x"c1",
  1879 => x"ca",
  1880 => x"f6",
  1881 => x"48",
  1882 => x"c1",
  1883 => x"78",
  1884 => x"c0",
  1885 => x"e4",
  1886 => x"87",
  1887 => x"c8",
  1888 => x"1e",
  1889 => x"c0",
  1890 => x"e7",
  1891 => x"f2",
  1892 => x"1e",
  1893 => x"c1",
  1894 => x"c3",
  1895 => x"e4",
  1896 => x"49",
  1897 => x"f9",
  1898 => x"f3",
  1899 => x"87",
  1900 => x"c8",
  1901 => x"86",
  1902 => x"70",
  1903 => x"98",
  1904 => x"02",
  1905 => x"c0",
  1906 => x"cf",
  1907 => x"87",
  1908 => x"c0",
  1909 => x"e5",
  1910 => x"f0",
  1911 => x"1e",
  1912 => x"c0",
  1913 => x"e2",
  1914 => x"ec",
  1915 => x"87",
  1916 => x"c4",
  1917 => x"86",
  1918 => x"c0",
  1919 => x"48",
  1920 => x"c6",
  1921 => x"cd",
  1922 => x"87",
  1923 => x"c1",
  1924 => x"ca",
  1925 => x"ec",
  1926 => x"97",
  1927 => x"bf",
  1928 => x"49",
  1929 => x"c1",
  1930 => x"d5",
  1931 => x"a9",
  1932 => x"05",
  1933 => x"c0",
  1934 => x"cd",
  1935 => x"87",
  1936 => x"c1",
  1937 => x"ca",
  1938 => x"ed",
  1939 => x"97",
  1940 => x"bf",
  1941 => x"49",
  1942 => x"c2",
  1943 => x"ea",
  1944 => x"a9",
  1945 => x"02",
  1946 => x"c0",
  1947 => x"c5",
  1948 => x"87",
  1949 => x"c0",
  1950 => x"48",
  1951 => x"c5",
  1952 => x"ee",
  1953 => x"87",
  1954 => x"c1",
  1955 => x"c2",
  1956 => x"ee",
  1957 => x"97",
  1958 => x"bf",
  1959 => x"49",
  1960 => x"c3",
  1961 => x"e9",
  1962 => x"a9",
  1963 => x"02",
  1964 => x"c0",
  1965 => x"d2",
  1966 => x"87",
  1967 => x"c1",
  1968 => x"c2",
  1969 => x"ee",
  1970 => x"97",
  1971 => x"bf",
  1972 => x"49",
  1973 => x"c3",
  1974 => x"eb",
  1975 => x"a9",
  1976 => x"02",
  1977 => x"c0",
  1978 => x"c5",
  1979 => x"87",
  1980 => x"c0",
  1981 => x"48",
  1982 => x"c5",
  1983 => x"cf",
  1984 => x"87",
  1985 => x"c1",
  1986 => x"c2",
  1987 => x"f9",
  1988 => x"97",
  1989 => x"bf",
  1990 => x"49",
  1991 => x"71",
  1992 => x"99",
  1993 => x"05",
  1994 => x"c0",
  1995 => x"cc",
  1996 => x"87",
  1997 => x"c1",
  1998 => x"c2",
  1999 => x"fa",
  2000 => x"97",
  2001 => x"bf",
  2002 => x"49",
  2003 => x"c2",
  2004 => x"a9",
  2005 => x"02",
  2006 => x"c0",
  2007 => x"c5",
  2008 => x"87",
  2009 => x"c0",
  2010 => x"48",
  2011 => x"c4",
  2012 => x"f2",
  2013 => x"87",
  2014 => x"c1",
  2015 => x"c2",
  2016 => x"fb",
  2017 => x"97",
  2018 => x"bf",
  2019 => x"48",
  2020 => x"c1",
  2021 => x"ca",
  2022 => x"f2",
  2023 => x"58",
  2024 => x"c1",
  2025 => x"ca",
  2026 => x"ee",
  2027 => x"bf",
  2028 => x"48",
  2029 => x"c1",
  2030 => x"88",
  2031 => x"c1",
  2032 => x"ca",
  2033 => x"f6",
  2034 => x"58",
  2035 => x"c1",
  2036 => x"c2",
  2037 => x"fc",
  2038 => x"97",
  2039 => x"bf",
  2040 => x"49",
  2041 => x"73",
  2042 => x"81",
  2043 => x"c1",
  2044 => x"c2",
  2045 => x"fd",
  2046 => x"97",
  2047 => x"bf",
  2048 => x"4a",
  2049 => x"c8",
  2050 => x"32",
  2051 => x"c1",
  2052 => x"cb",
  2053 => x"c2",
  2054 => x"48",
  2055 => x"72",
  2056 => x"a1",
  2057 => x"78",
  2058 => x"c1",
  2059 => x"c2",
  2060 => x"fe",
  2061 => x"97",
  2062 => x"bf",
  2063 => x"48",
  2064 => x"c1",
  2065 => x"cb",
  2066 => x"da",
  2067 => x"58",
  2068 => x"c1",
  2069 => x"ca",
  2070 => x"f6",
  2071 => x"bf",
  2072 => x"02",
  2073 => x"c2",
  2074 => x"e2",
  2075 => x"87",
  2076 => x"c8",
  2077 => x"1e",
  2078 => x"c0",
  2079 => x"e6",
  2080 => x"cd",
  2081 => x"1e",
  2082 => x"c1",
  2083 => x"c4",
  2084 => x"c0",
  2085 => x"49",
  2086 => x"f6",
  2087 => x"f6",
  2088 => x"87",
  2089 => x"c8",
  2090 => x"86",
  2091 => x"70",
  2092 => x"98",
  2093 => x"02",
  2094 => x"c0",
  2095 => x"c5",
  2096 => x"87",
  2097 => x"c0",
  2098 => x"48",
  2099 => x"c3",
  2100 => x"da",
  2101 => x"87",
  2102 => x"c1",
  2103 => x"ca",
  2104 => x"ee",
  2105 => x"bf",
  2106 => x"48",
  2107 => x"c4",
  2108 => x"30",
  2109 => x"c1",
  2110 => x"cb",
  2111 => x"de",
  2112 => x"58",
  2113 => x"c1",
  2114 => x"ca",
  2115 => x"ee",
  2116 => x"bf",
  2117 => x"4a",
  2118 => x"c1",
  2119 => x"cb",
  2120 => x"d6",
  2121 => x"5a",
  2122 => x"c1",
  2123 => x"c3",
  2124 => x"d3",
  2125 => x"97",
  2126 => x"bf",
  2127 => x"49",
  2128 => x"c8",
  2129 => x"31",
  2130 => x"c1",
  2131 => x"c3",
  2132 => x"d2",
  2133 => x"97",
  2134 => x"bf",
  2135 => x"4b",
  2136 => x"73",
  2137 => x"a1",
  2138 => x"49",
  2139 => x"c1",
  2140 => x"c3",
  2141 => x"d4",
  2142 => x"97",
  2143 => x"bf",
  2144 => x"4b",
  2145 => x"d0",
  2146 => x"33",
  2147 => x"73",
  2148 => x"a1",
  2149 => x"49",
  2150 => x"c1",
  2151 => x"c3",
  2152 => x"d5",
  2153 => x"97",
  2154 => x"bf",
  2155 => x"4b",
  2156 => x"d8",
  2157 => x"33",
  2158 => x"73",
  2159 => x"a1",
  2160 => x"49",
  2161 => x"c1",
  2162 => x"cb",
  2163 => x"e2",
  2164 => x"59",
  2165 => x"c1",
  2166 => x"cb",
  2167 => x"d6",
  2168 => x"bf",
  2169 => x"91",
  2170 => x"c1",
  2171 => x"cb",
  2172 => x"c2",
  2173 => x"bf",
  2174 => x"81",
  2175 => x"c1",
  2176 => x"cb",
  2177 => x"ca",
  2178 => x"59",
  2179 => x"c1",
  2180 => x"c3",
  2181 => x"db",
  2182 => x"97",
  2183 => x"bf",
  2184 => x"4b",
  2185 => x"c8",
  2186 => x"33",
  2187 => x"c1",
  2188 => x"c3",
  2189 => x"da",
  2190 => x"97",
  2191 => x"bf",
  2192 => x"4c",
  2193 => x"74",
  2194 => x"a3",
  2195 => x"4b",
  2196 => x"c1",
  2197 => x"c3",
  2198 => x"dc",
  2199 => x"97",
  2200 => x"bf",
  2201 => x"4c",
  2202 => x"d0",
  2203 => x"34",
  2204 => x"74",
  2205 => x"a3",
  2206 => x"4b",
  2207 => x"c1",
  2208 => x"c3",
  2209 => x"dd",
  2210 => x"97",
  2211 => x"bf",
  2212 => x"4c",
  2213 => x"cf",
  2214 => x"9c",
  2215 => x"d8",
  2216 => x"34",
  2217 => x"74",
  2218 => x"a3",
  2219 => x"4b",
  2220 => x"c1",
  2221 => x"cb",
  2222 => x"ce",
  2223 => x"5b",
  2224 => x"c2",
  2225 => x"8b",
  2226 => x"73",
  2227 => x"92",
  2228 => x"c1",
  2229 => x"cb",
  2230 => x"ce",
  2231 => x"48",
  2232 => x"72",
  2233 => x"a1",
  2234 => x"78",
  2235 => x"c1",
  2236 => x"d0",
  2237 => x"87",
  2238 => x"c1",
  2239 => x"c3",
  2240 => x"c0",
  2241 => x"97",
  2242 => x"bf",
  2243 => x"49",
  2244 => x"c8",
  2245 => x"31",
  2246 => x"c1",
  2247 => x"c2",
  2248 => x"ff",
  2249 => x"97",
  2250 => x"bf",
  2251 => x"4a",
  2252 => x"72",
  2253 => x"a1",
  2254 => x"49",
  2255 => x"c1",
  2256 => x"cb",
  2257 => x"de",
  2258 => x"59",
  2259 => x"c5",
  2260 => x"31",
  2261 => x"c7",
  2262 => x"ff",
  2263 => x"81",
  2264 => x"c9",
  2265 => x"29",
  2266 => x"c1",
  2267 => x"cb",
  2268 => x"d6",
  2269 => x"59",
  2270 => x"c1",
  2271 => x"c3",
  2272 => x"c5",
  2273 => x"97",
  2274 => x"bf",
  2275 => x"4a",
  2276 => x"c8",
  2277 => x"32",
  2278 => x"c1",
  2279 => x"c3",
  2280 => x"c4",
  2281 => x"97",
  2282 => x"bf",
  2283 => x"4b",
  2284 => x"73",
  2285 => x"a2",
  2286 => x"4a",
  2287 => x"c1",
  2288 => x"cb",
  2289 => x"e2",
  2290 => x"5a",
  2291 => x"c1",
  2292 => x"cb",
  2293 => x"d6",
  2294 => x"bf",
  2295 => x"92",
  2296 => x"c1",
  2297 => x"cb",
  2298 => x"c2",
  2299 => x"bf",
  2300 => x"82",
  2301 => x"c1",
  2302 => x"cb",
  2303 => x"d2",
  2304 => x"5a",
  2305 => x"c1",
  2306 => x"cb",
  2307 => x"ca",
  2308 => x"48",
  2309 => x"c0",
  2310 => x"78",
  2311 => x"c1",
  2312 => x"cb",
  2313 => x"c6",
  2314 => x"48",
  2315 => x"72",
  2316 => x"a1",
  2317 => x"78",
  2318 => x"c1",
  2319 => x"48",
  2320 => x"f4",
  2321 => x"c6",
  2322 => x"87",
  2323 => x"4e",
  2324 => x"6f",
  2325 => x"20",
  2326 => x"70",
  2327 => x"61",
  2328 => x"72",
  2329 => x"74",
  2330 => x"69",
  2331 => x"74",
  2332 => x"69",
  2333 => x"6f",
  2334 => x"6e",
  2335 => x"20",
  2336 => x"73",
  2337 => x"69",
  2338 => x"67",
  2339 => x"6e",
  2340 => x"61",
  2341 => x"74",
  2342 => x"75",
  2343 => x"72",
  2344 => x"65",
  2345 => x"20",
  2346 => x"66",
  2347 => x"6f",
  2348 => x"75",
  2349 => x"6e",
  2350 => x"64",
  2351 => x"0a",
  2352 => x"00",
  2353 => x"52",
  2354 => x"65",
  2355 => x"61",
  2356 => x"64",
  2357 => x"69",
  2358 => x"6e",
  2359 => x"67",
  2360 => x"20",
  2361 => x"62",
  2362 => x"6f",
  2363 => x"6f",
  2364 => x"74",
  2365 => x"20",
  2366 => x"73",
  2367 => x"65",
  2368 => x"63",
  2369 => x"74",
  2370 => x"6f",
  2371 => x"72",
  2372 => x"20",
  2373 => x"25",
  2374 => x"64",
  2375 => x"0a",
  2376 => x"00",
  2377 => x"52",
  2378 => x"65",
  2379 => x"61",
  2380 => x"64",
  2381 => x"20",
  2382 => x"62",
  2383 => x"6f",
  2384 => x"6f",
  2385 => x"74",
  2386 => x"20",
  2387 => x"73",
  2388 => x"65",
  2389 => x"63",
  2390 => x"74",
  2391 => x"6f",
  2392 => x"72",
  2393 => x"20",
  2394 => x"66",
  2395 => x"72",
  2396 => x"6f",
  2397 => x"6d",
  2398 => x"20",
  2399 => x"66",
  2400 => x"69",
  2401 => x"72",
  2402 => x"73",
  2403 => x"74",
  2404 => x"20",
  2405 => x"70",
  2406 => x"61",
  2407 => x"72",
  2408 => x"74",
  2409 => x"69",
  2410 => x"74",
  2411 => x"69",
  2412 => x"6f",
  2413 => x"6e",
  2414 => x"0a",
  2415 => x"00",
  2416 => x"55",
  2417 => x"6e",
  2418 => x"73",
  2419 => x"75",
  2420 => x"70",
  2421 => x"70",
  2422 => x"6f",
  2423 => x"72",
  2424 => x"74",
  2425 => x"65",
  2426 => x"64",
  2427 => x"20",
  2428 => x"70",
  2429 => x"61",
  2430 => x"72",
  2431 => x"74",
  2432 => x"69",
  2433 => x"74",
  2434 => x"69",
  2435 => x"6f",
  2436 => x"6e",
  2437 => x"20",
  2438 => x"74",
  2439 => x"79",
  2440 => x"70",
  2441 => x"65",
  2442 => x"21",
  2443 => x"0d",
  2444 => x"00",
  2445 => x"46",
  2446 => x"41",
  2447 => x"54",
  2448 => x"33",
  2449 => x"32",
  2450 => x"20",
  2451 => x"20",
  2452 => x"20",
  2453 => x"00",
  2454 => x"52",
  2455 => x"65",
  2456 => x"61",
  2457 => x"64",
  2458 => x"69",
  2459 => x"6e",
  2460 => x"67",
  2461 => x"20",
  2462 => x"4d",
  2463 => x"42",
  2464 => x"52",
  2465 => x"0a",
  2466 => x"00",
  2467 => x"46",
  2468 => x"41",
  2469 => x"54",
  2470 => x"31",
  2471 => x"36",
  2472 => x"20",
  2473 => x"20",
  2474 => x"20",
  2475 => x"00",
  2476 => x"46",
  2477 => x"41",
  2478 => x"54",
  2479 => x"33",
  2480 => x"32",
  2481 => x"20",
  2482 => x"20",
  2483 => x"20",
  2484 => x"00",
  2485 => x"46",
  2486 => x"41",
  2487 => x"54",
  2488 => x"31",
  2489 => x"32",
  2490 => x"20",
  2491 => x"20",
  2492 => x"20",
  2493 => x"00",
  2494 => x"50",
  2495 => x"61",
  2496 => x"72",
  2497 => x"74",
  2498 => x"69",
  2499 => x"74",
  2500 => x"69",
  2501 => x"6f",
  2502 => x"6e",
  2503 => x"63",
  2504 => x"6f",
  2505 => x"75",
  2506 => x"6e",
  2507 => x"74",
  2508 => x"20",
  2509 => x"25",
  2510 => x"64",
  2511 => x"0a",
  2512 => x"00",
  2513 => x"48",
  2514 => x"75",
  2515 => x"6e",
  2516 => x"74",
  2517 => x"69",
  2518 => x"6e",
  2519 => x"67",
  2520 => x"20",
  2521 => x"66",
  2522 => x"6f",
  2523 => x"72",
  2524 => x"20",
  2525 => x"66",
  2526 => x"69",
  2527 => x"6c",
  2528 => x"65",
  2529 => x"73",
  2530 => x"79",
  2531 => x"73",
  2532 => x"74",
  2533 => x"65",
  2534 => x"6d",
  2535 => x"0a",
  2536 => x"00",
  2537 => x"46",
  2538 => x"41",
  2539 => x"54",
  2540 => x"33",
  2541 => x"32",
  2542 => x"20",
  2543 => x"20",
  2544 => x"20",
  2545 => x"00",
  2546 => x"46",
  2547 => x"41",
  2548 => x"54",
  2549 => x"31",
  2550 => x"36",
  2551 => x"20",
  2552 => x"20",
  2553 => x"20",
  2554 => x"00",
  2555 => x"52",
  2556 => x"65",
  2557 => x"61",
  2558 => x"64",
  2559 => x"69",
  2560 => x"6e",
  2561 => x"67",
  2562 => x"20",
  2563 => x"64",
  2564 => x"69",
  2565 => x"72",
  2566 => x"65",
  2567 => x"63",
  2568 => x"74",
  2569 => x"6f",
  2570 => x"72",
  2571 => x"79",
  2572 => x"20",
  2573 => x"73",
  2574 => x"65",
  2575 => x"63",
  2576 => x"74",
  2577 => x"6f",
  2578 => x"72",
  2579 => x"20",
  2580 => x"25",
  2581 => x"64",
  2582 => x"0a",
  2583 => x"00",
  2584 => x"66",
  2585 => x"69",
  2586 => x"6c",
  2587 => x"65",
  2588 => x"20",
  2589 => x"22",
  2590 => x"25",
  2591 => x"73",
  2592 => x"22",
  2593 => x"20",
  2594 => x"66",
  2595 => x"6f",
  2596 => x"75",
  2597 => x"6e",
  2598 => x"64",
  2599 => x"0d",
  2600 => x"00",
  2601 => x"47",
  2602 => x"65",
  2603 => x"74",
  2604 => x"46",
  2605 => x"41",
  2606 => x"54",
  2607 => x"4c",
  2608 => x"69",
  2609 => x"6e",
  2610 => x"6b",
  2611 => x"20",
  2612 => x"72",
  2613 => x"65",
  2614 => x"74",
  2615 => x"75",
  2616 => x"72",
  2617 => x"6e",
  2618 => x"65",
  2619 => x"64",
  2620 => x"20",
  2621 => x"25",
  2622 => x"64",
  2623 => x"0a",
  2624 => x"00",
  2625 => x"43",
  2626 => x"61",
  2627 => x"6e",
  2628 => x"27",
  2629 => x"74",
  2630 => x"20",
  2631 => x"6f",
  2632 => x"70",
  2633 => x"65",
  2634 => x"6e",
  2635 => x"20",
  2636 => x"25",
  2637 => x"73",
  2638 => x"0a",
  2639 => x"00",
  2640 => x"0e",
  2641 => x"5e",
  2642 => x"5b",
  2643 => x"5c",
  2644 => x"5d",
  2645 => x"0e",
  2646 => x"71",
  2647 => x"4a",
  2648 => x"c1",
  2649 => x"ca",
  2650 => x"f6",
  2651 => x"bf",
  2652 => x"02",
  2653 => x"cc",
  2654 => x"87",
  2655 => x"72",
  2656 => x"4b",
  2657 => x"c7",
  2658 => x"b7",
  2659 => x"2b",
  2660 => x"72",
  2661 => x"4c",
  2662 => x"c1",
  2663 => x"ff",
  2664 => x"9c",
  2665 => x"ca",
  2666 => x"87",
  2667 => x"72",
  2668 => x"4b",
  2669 => x"c8",
  2670 => x"b7",
  2671 => x"2b",
  2672 => x"72",
  2673 => x"4c",
  2674 => x"c3",
  2675 => x"ff",
  2676 => x"9c",
  2677 => x"c1",
  2678 => x"cb",
  2679 => x"e6",
  2680 => x"bf",
  2681 => x"ab",
  2682 => x"02",
  2683 => x"de",
  2684 => x"87",
  2685 => x"c1",
  2686 => x"c2",
  2687 => x"ee",
  2688 => x"1e",
  2689 => x"c1",
  2690 => x"cb",
  2691 => x"c2",
  2692 => x"bf",
  2693 => x"49",
  2694 => x"73",
  2695 => x"81",
  2696 => x"ea",
  2697 => x"c1",
  2698 => x"87",
  2699 => x"c4",
  2700 => x"86",
  2701 => x"70",
  2702 => x"98",
  2703 => x"05",
  2704 => x"c5",
  2705 => x"87",
  2706 => x"c0",
  2707 => x"48",
  2708 => x"c0",
  2709 => x"f6",
  2710 => x"87",
  2711 => x"c1",
  2712 => x"cb",
  2713 => x"ea",
  2714 => x"5b",
  2715 => x"c1",
  2716 => x"ca",
  2717 => x"f6",
  2718 => x"bf",
  2719 => x"02",
  2720 => x"d9",
  2721 => x"87",
  2722 => x"74",
  2723 => x"4a",
  2724 => x"c4",
  2725 => x"92",
  2726 => x"c1",
  2727 => x"c2",
  2728 => x"ee",
  2729 => x"82",
  2730 => x"6a",
  2731 => x"49",
  2732 => x"eb",
  2733 => x"dc",
  2734 => x"87",
  2735 => x"70",
  2736 => x"49",
  2737 => x"71",
  2738 => x"4d",
  2739 => x"cf",
  2740 => x"ff",
  2741 => x"ff",
  2742 => x"ff",
  2743 => x"ff",
  2744 => x"9d",
  2745 => x"d0",
  2746 => x"87",
  2747 => x"74",
  2748 => x"4a",
  2749 => x"c2",
  2750 => x"92",
  2751 => x"c1",
  2752 => x"c2",
  2753 => x"ee",
  2754 => x"82",
  2755 => x"9f",
  2756 => x"6a",
  2757 => x"49",
  2758 => x"eb",
  2759 => x"fc",
  2760 => x"87",
  2761 => x"70",
  2762 => x"4d",
  2763 => x"75",
  2764 => x"48",
  2765 => x"ed",
  2766 => x"c9",
  2767 => x"87",
  2768 => x"0e",
  2769 => x"5e",
  2770 => x"5b",
  2771 => x"5c",
  2772 => x"5d",
  2773 => x"0e",
  2774 => x"f4",
  2775 => x"86",
  2776 => x"71",
  2777 => x"4c",
  2778 => x"c0",
  2779 => x"4b",
  2780 => x"c1",
  2781 => x"cb",
  2782 => x"e6",
  2783 => x"48",
  2784 => x"ff",
  2785 => x"78",
  2786 => x"c1",
  2787 => x"cb",
  2788 => x"ca",
  2789 => x"bf",
  2790 => x"4d",
  2791 => x"c1",
  2792 => x"cb",
  2793 => x"ce",
  2794 => x"bf",
  2795 => x"7e",
  2796 => x"c1",
  2797 => x"ca",
  2798 => x"f6",
  2799 => x"bf",
  2800 => x"02",
  2801 => x"c9",
  2802 => x"87",
  2803 => x"c1",
  2804 => x"ca",
  2805 => x"ee",
  2806 => x"bf",
  2807 => x"4a",
  2808 => x"c4",
  2809 => x"32",
  2810 => x"c7",
  2811 => x"87",
  2812 => x"c1",
  2813 => x"cb",
  2814 => x"d2",
  2815 => x"bf",
  2816 => x"4a",
  2817 => x"c4",
  2818 => x"32",
  2819 => x"c8",
  2820 => x"a6",
  2821 => x"5a",
  2822 => x"c8",
  2823 => x"a6",
  2824 => x"48",
  2825 => x"c0",
  2826 => x"78",
  2827 => x"c4",
  2828 => x"66",
  2829 => x"48",
  2830 => x"c0",
  2831 => x"a8",
  2832 => x"06",
  2833 => x"c3",
  2834 => x"cf",
  2835 => x"87",
  2836 => x"c8",
  2837 => x"66",
  2838 => x"49",
  2839 => x"cf",
  2840 => x"99",
  2841 => x"05",
  2842 => x"c0",
  2843 => x"e3",
  2844 => x"87",
  2845 => x"6e",
  2846 => x"1e",
  2847 => x"c0",
  2848 => x"e7",
  2849 => x"fb",
  2850 => x"1e",
  2851 => x"d4",
  2852 => x"c2",
  2853 => x"87",
  2854 => x"c1",
  2855 => x"c2",
  2856 => x"ee",
  2857 => x"1e",
  2858 => x"cc",
  2859 => x"66",
  2860 => x"49",
  2861 => x"48",
  2862 => x"c1",
  2863 => x"80",
  2864 => x"d0",
  2865 => x"a6",
  2866 => x"58",
  2867 => x"71",
  2868 => x"49",
  2869 => x"e7",
  2870 => x"d4",
  2871 => x"87",
  2872 => x"cc",
  2873 => x"86",
  2874 => x"c1",
  2875 => x"c2",
  2876 => x"ee",
  2877 => x"4b",
  2878 => x"c3",
  2879 => x"87",
  2880 => x"c0",
  2881 => x"e0",
  2882 => x"83",
  2883 => x"97",
  2884 => x"6b",
  2885 => x"49",
  2886 => x"71",
  2887 => x"99",
  2888 => x"02",
  2889 => x"c2",
  2890 => x"c5",
  2891 => x"87",
  2892 => x"97",
  2893 => x"6b",
  2894 => x"49",
  2895 => x"c3",
  2896 => x"e5",
  2897 => x"a9",
  2898 => x"02",
  2899 => x"c1",
  2900 => x"fb",
  2901 => x"87",
  2902 => x"cb",
  2903 => x"a3",
  2904 => x"49",
  2905 => x"97",
  2906 => x"69",
  2907 => x"49",
  2908 => x"d8",
  2909 => x"99",
  2910 => x"05",
  2911 => x"c1",
  2912 => x"ef",
  2913 => x"87",
  2914 => x"cb",
  2915 => x"1e",
  2916 => x"c0",
  2917 => x"e0",
  2918 => x"66",
  2919 => x"1e",
  2920 => x"73",
  2921 => x"49",
  2922 => x"e9",
  2923 => x"f2",
  2924 => x"87",
  2925 => x"c8",
  2926 => x"86",
  2927 => x"70",
  2928 => x"98",
  2929 => x"05",
  2930 => x"c1",
  2931 => x"dc",
  2932 => x"87",
  2933 => x"dc",
  2934 => x"a3",
  2935 => x"4a",
  2936 => x"6a",
  2937 => x"49",
  2938 => x"e8",
  2939 => x"ce",
  2940 => x"87",
  2941 => x"70",
  2942 => x"4a",
  2943 => x"c4",
  2944 => x"a4",
  2945 => x"49",
  2946 => x"72",
  2947 => x"79",
  2948 => x"da",
  2949 => x"a3",
  2950 => x"4a",
  2951 => x"9f",
  2952 => x"6a",
  2953 => x"49",
  2954 => x"e8",
  2955 => x"f8",
  2956 => x"87",
  2957 => x"c4",
  2958 => x"a6",
  2959 => x"58",
  2960 => x"c1",
  2961 => x"ca",
  2962 => x"f6",
  2963 => x"bf",
  2964 => x"02",
  2965 => x"d8",
  2966 => x"87",
  2967 => x"d4",
  2968 => x"a3",
  2969 => x"4a",
  2970 => x"9f",
  2971 => x"6a",
  2972 => x"49",
  2973 => x"e8",
  2974 => x"e5",
  2975 => x"87",
  2976 => x"70",
  2977 => x"49",
  2978 => x"c0",
  2979 => x"ff",
  2980 => x"ff",
  2981 => x"99",
  2982 => x"71",
  2983 => x"48",
  2984 => x"d0",
  2985 => x"30",
  2986 => x"c8",
  2987 => x"a6",
  2988 => x"58",
  2989 => x"c5",
  2990 => x"87",
  2991 => x"c4",
  2992 => x"a6",
  2993 => x"48",
  2994 => x"c0",
  2995 => x"78",
  2996 => x"c4",
  2997 => x"66",
  2998 => x"4a",
  2999 => x"6e",
  3000 => x"82",
  3001 => x"c8",
  3002 => x"a4",
  3003 => x"49",
  3004 => x"72",
  3005 => x"79",
  3006 => x"c0",
  3007 => x"7c",
  3008 => x"dc",
  3009 => x"66",
  3010 => x"1e",
  3011 => x"c0",
  3012 => x"e8",
  3013 => x"d8",
  3014 => x"1e",
  3015 => x"d1",
  3016 => x"de",
  3017 => x"87",
  3018 => x"c8",
  3019 => x"86",
  3020 => x"c1",
  3021 => x"48",
  3022 => x"c1",
  3023 => x"d0",
  3024 => x"87",
  3025 => x"c8",
  3026 => x"66",
  3027 => x"48",
  3028 => x"c1",
  3029 => x"80",
  3030 => x"cc",
  3031 => x"a6",
  3032 => x"58",
  3033 => x"c8",
  3034 => x"66",
  3035 => x"48",
  3036 => x"c4",
  3037 => x"66",
  3038 => x"a8",
  3039 => x"04",
  3040 => x"fc",
  3041 => x"f1",
  3042 => x"87",
  3043 => x"c1",
  3044 => x"ca",
  3045 => x"f6",
  3046 => x"bf",
  3047 => x"02",
  3048 => x"c0",
  3049 => x"f4",
  3050 => x"87",
  3051 => x"75",
  3052 => x"49",
  3053 => x"f9",
  3054 => x"e0",
  3055 => x"87",
  3056 => x"70",
  3057 => x"4d",
  3058 => x"75",
  3059 => x"1e",
  3060 => x"c0",
  3061 => x"e8",
  3062 => x"e9",
  3063 => x"1e",
  3064 => x"d0",
  3065 => x"ed",
  3066 => x"87",
  3067 => x"c8",
  3068 => x"86",
  3069 => x"75",
  3070 => x"49",
  3071 => x"cf",
  3072 => x"ff",
  3073 => x"ff",
  3074 => x"ff",
  3075 => x"f8",
  3076 => x"99",
  3077 => x"a9",
  3078 => x"02",
  3079 => x"d6",
  3080 => x"87",
  3081 => x"75",
  3082 => x"49",
  3083 => x"c2",
  3084 => x"89",
  3085 => x"c1",
  3086 => x"ca",
  3087 => x"ee",
  3088 => x"bf",
  3089 => x"91",
  3090 => x"c1",
  3091 => x"cb",
  3092 => x"c6",
  3093 => x"bf",
  3094 => x"48",
  3095 => x"71",
  3096 => x"80",
  3097 => x"c4",
  3098 => x"a6",
  3099 => x"58",
  3100 => x"fb",
  3101 => x"e7",
  3102 => x"87",
  3103 => x"c0",
  3104 => x"48",
  3105 => x"f4",
  3106 => x"8e",
  3107 => x"e7",
  3108 => x"f3",
  3109 => x"87",
  3110 => x"0e",
  3111 => x"5e",
  3112 => x"5b",
  3113 => x"5c",
  3114 => x"5d",
  3115 => x"0e",
  3116 => x"1e",
  3117 => x"71",
  3118 => x"4b",
  3119 => x"73",
  3120 => x"1e",
  3121 => x"c1",
  3122 => x"cb",
  3123 => x"ea",
  3124 => x"49",
  3125 => x"fa",
  3126 => x"d8",
  3127 => x"87",
  3128 => x"c4",
  3129 => x"86",
  3130 => x"70",
  3131 => x"98",
  3132 => x"02",
  3133 => x"c1",
  3134 => x"f7",
  3135 => x"87",
  3136 => x"c1",
  3137 => x"cb",
  3138 => x"ee",
  3139 => x"bf",
  3140 => x"49",
  3141 => x"c7",
  3142 => x"ff",
  3143 => x"81",
  3144 => x"c9",
  3145 => x"29",
  3146 => x"c4",
  3147 => x"a6",
  3148 => x"59",
  3149 => x"c0",
  3150 => x"4d",
  3151 => x"4c",
  3152 => x"6e",
  3153 => x"48",
  3154 => x"c0",
  3155 => x"b7",
  3156 => x"a8",
  3157 => x"06",
  3158 => x"c1",
  3159 => x"ed",
  3160 => x"87",
  3161 => x"c1",
  3162 => x"cb",
  3163 => x"c6",
  3164 => x"bf",
  3165 => x"49",
  3166 => x"c1",
  3167 => x"cb",
  3168 => x"f2",
  3169 => x"bf",
  3170 => x"4a",
  3171 => x"c2",
  3172 => x"8a",
  3173 => x"c1",
  3174 => x"ca",
  3175 => x"ee",
  3176 => x"bf",
  3177 => x"92",
  3178 => x"72",
  3179 => x"a1",
  3180 => x"49",
  3181 => x"c1",
  3182 => x"ca",
  3183 => x"f2",
  3184 => x"bf",
  3185 => x"4a",
  3186 => x"74",
  3187 => x"9a",
  3188 => x"72",
  3189 => x"a1",
  3190 => x"49",
  3191 => x"d4",
  3192 => x"66",
  3193 => x"1e",
  3194 => x"71",
  3195 => x"49",
  3196 => x"e2",
  3197 => x"cd",
  3198 => x"87",
  3199 => x"c4",
  3200 => x"86",
  3201 => x"70",
  3202 => x"98",
  3203 => x"05",
  3204 => x"c5",
  3205 => x"87",
  3206 => x"c0",
  3207 => x"48",
  3208 => x"c1",
  3209 => x"c0",
  3210 => x"87",
  3211 => x"c1",
  3212 => x"84",
  3213 => x"c1",
  3214 => x"ca",
  3215 => x"f2",
  3216 => x"bf",
  3217 => x"49",
  3218 => x"74",
  3219 => x"99",
  3220 => x"05",
  3221 => x"cc",
  3222 => x"87",
  3223 => x"c1",
  3224 => x"cb",
  3225 => x"f2",
  3226 => x"bf",
  3227 => x"49",
  3228 => x"f6",
  3229 => x"f1",
  3230 => x"87",
  3231 => x"c1",
  3232 => x"cb",
  3233 => x"f6",
  3234 => x"58",
  3235 => x"d4",
  3236 => x"66",
  3237 => x"48",
  3238 => x"c8",
  3239 => x"c0",
  3240 => x"80",
  3241 => x"d8",
  3242 => x"a6",
  3243 => x"58",
  3244 => x"c1",
  3245 => x"85",
  3246 => x"6e",
  3247 => x"b7",
  3248 => x"ad",
  3249 => x"04",
  3250 => x"fe",
  3251 => x"e4",
  3252 => x"87",
  3253 => x"cf",
  3254 => x"87",
  3255 => x"73",
  3256 => x"1e",
  3257 => x"c0",
  3258 => x"e9",
  3259 => x"c1",
  3260 => x"1e",
  3261 => x"cd",
  3262 => x"e8",
  3263 => x"87",
  3264 => x"c8",
  3265 => x"86",
  3266 => x"c0",
  3267 => x"48",
  3268 => x"c5",
  3269 => x"87",
  3270 => x"c1",
  3271 => x"cb",
  3272 => x"ee",
  3273 => x"bf",
  3274 => x"48",
  3275 => x"26",
  3276 => x"e5",
  3277 => x"ca",
  3278 => x"87",
  3279 => x"1e",
  3280 => x"f1",
  3281 => x"09",
  3282 => x"97",
  3283 => x"79",
  3284 => x"09",
  3285 => x"71",
  3286 => x"48",
  3287 => x"26",
  3288 => x"4f",
  3289 => x"0e",
  3290 => x"5e",
  3291 => x"5b",
  3292 => x"5c",
  3293 => x"0e",
  3294 => x"71",
  3295 => x"4b",
  3296 => x"c0",
  3297 => x"4c",
  3298 => x"13",
  3299 => x"4a",
  3300 => x"72",
  3301 => x"9a",
  3302 => x"02",
  3303 => x"cd",
  3304 => x"87",
  3305 => x"72",
  3306 => x"49",
  3307 => x"e2",
  3308 => x"87",
  3309 => x"c1",
  3310 => x"84",
  3311 => x"13",
  3312 => x"4a",
  3313 => x"72",
  3314 => x"9a",
  3315 => x"05",
  3316 => x"f3",
  3317 => x"87",
  3318 => x"74",
  3319 => x"48",
  3320 => x"c2",
  3321 => x"87",
  3322 => x"26",
  3323 => x"4d",
  3324 => x"26",
  3325 => x"4c",
  3326 => x"26",
  3327 => x"4b",
  3328 => x"26",
  3329 => x"4f",
  3330 => x"0e",
  3331 => x"5e",
  3332 => x"5b",
  3333 => x"5c",
  3334 => x"5d",
  3335 => x"0e",
  3336 => x"71",
  3337 => x"4b",
  3338 => x"73",
  3339 => x"4c",
  3340 => x"d0",
  3341 => x"66",
  3342 => x"48",
  3343 => x"c2",
  3344 => x"28",
  3345 => x"d4",
  3346 => x"a6",
  3347 => x"58",
  3348 => x"d0",
  3349 => x"66",
  3350 => x"49",
  3351 => x"48",
  3352 => x"c1",
  3353 => x"88",
  3354 => x"d4",
  3355 => x"a6",
  3356 => x"58",
  3357 => x"71",
  3358 => x"99",
  3359 => x"02",
  3360 => x"c1",
  3361 => x"c4",
  3362 => x"87",
  3363 => x"24",
  3364 => x"4d",
  3365 => x"c0",
  3366 => x"4b",
  3367 => x"75",
  3368 => x"4a",
  3369 => x"dc",
  3370 => x"2a",
  3371 => x"c0",
  3372 => x"f0",
  3373 => x"82",
  3374 => x"c0",
  3375 => x"f9",
  3376 => x"aa",
  3377 => x"06",
  3378 => x"c2",
  3379 => x"87",
  3380 => x"c7",
  3381 => x"82",
  3382 => x"72",
  3383 => x"49",
  3384 => x"fe",
  3385 => x"d4",
  3386 => x"87",
  3387 => x"c4",
  3388 => x"35",
  3389 => x"c1",
  3390 => x"83",
  3391 => x"c8",
  3392 => x"b7",
  3393 => x"ab",
  3394 => x"04",
  3395 => x"e2",
  3396 => x"87",
  3397 => x"c0",
  3398 => x"e0",
  3399 => x"49",
  3400 => x"fe",
  3401 => x"c4",
  3402 => x"87",
  3403 => x"d0",
  3404 => x"66",
  3405 => x"49",
  3406 => x"c3",
  3407 => x"99",
  3408 => x"05",
  3409 => x"c5",
  3410 => x"87",
  3411 => x"ca",
  3412 => x"49",
  3413 => x"fd",
  3414 => x"f7",
  3415 => x"87",
  3416 => x"d0",
  3417 => x"66",
  3418 => x"49",
  3419 => x"48",
  3420 => x"c1",
  3421 => x"88",
  3422 => x"d4",
  3423 => x"a6",
  3424 => x"58",
  3425 => x"71",
  3426 => x"99",
  3427 => x"05",
  3428 => x"fe",
  3429 => x"fc",
  3430 => x"87",
  3431 => x"ca",
  3432 => x"49",
  3433 => x"fd",
  3434 => x"e3",
  3435 => x"87",
  3436 => x"26",
  3437 => x"4d",
  3438 => x"26",
  3439 => x"4c",
  3440 => x"26",
  3441 => x"4b",
  3442 => x"26",
  3443 => x"4f",
  3444 => x"0e",
  3445 => x"5e",
  3446 => x"5b",
  3447 => x"5c",
  3448 => x"5d",
  3449 => x"0e",
  3450 => x"fc",
  3451 => x"86",
  3452 => x"71",
  3453 => x"4a",
  3454 => x"c0",
  3455 => x"e0",
  3456 => x"66",
  3457 => x"4c",
  3458 => x"c1",
  3459 => x"cb",
  3460 => x"f6",
  3461 => x"4b",
  3462 => x"c0",
  3463 => x"7e",
  3464 => x"72",
  3465 => x"9a",
  3466 => x"05",
  3467 => x"ce",
  3468 => x"87",
  3469 => x"c1",
  3470 => x"cb",
  3471 => x"f7",
  3472 => x"4b",
  3473 => x"c1",
  3474 => x"cb",
  3475 => x"f6",
  3476 => x"48",
  3477 => x"c0",
  3478 => x"f0",
  3479 => x"50",
  3480 => x"c1",
  3481 => x"d2",
  3482 => x"87",
  3483 => x"72",
  3484 => x"9a",
  3485 => x"02",
  3486 => x"c0",
  3487 => x"e9",
  3488 => x"87",
  3489 => x"d4",
  3490 => x"66",
  3491 => x"4d",
  3492 => x"72",
  3493 => x"1e",
  3494 => x"72",
  3495 => x"49",
  3496 => x"75",
  3497 => x"4a",
  3498 => x"ca",
  3499 => x"cf",
  3500 => x"87",
  3501 => x"26",
  3502 => x"4a",
  3503 => x"c0",
  3504 => x"f8",
  3505 => x"de",
  3506 => x"81",
  3507 => x"11",
  3508 => x"53",
  3509 => x"71",
  3510 => x"1e",
  3511 => x"72",
  3512 => x"49",
  3513 => x"75",
  3514 => x"4a",
  3515 => x"c9",
  3516 => x"fe",
  3517 => x"87",
  3518 => x"70",
  3519 => x"4a",
  3520 => x"26",
  3521 => x"49",
  3522 => x"c1",
  3523 => x"8c",
  3524 => x"72",
  3525 => x"9a",
  3526 => x"05",
  3527 => x"ff",
  3528 => x"da",
  3529 => x"87",
  3530 => x"c0",
  3531 => x"b7",
  3532 => x"ac",
  3533 => x"06",
  3534 => x"dd",
  3535 => x"87",
  3536 => x"c0",
  3537 => x"e4",
  3538 => x"66",
  3539 => x"02",
  3540 => x"c5",
  3541 => x"87",
  3542 => x"c0",
  3543 => x"f0",
  3544 => x"4a",
  3545 => x"c3",
  3546 => x"87",
  3547 => x"c0",
  3548 => x"e0",
  3549 => x"4a",
  3550 => x"73",
  3551 => x"0a",
  3552 => x"97",
  3553 => x"7a",
  3554 => x"0a",
  3555 => x"c1",
  3556 => x"83",
  3557 => x"8c",
  3558 => x"c0",
  3559 => x"b7",
  3560 => x"ac",
  3561 => x"01",
  3562 => x"ff",
  3563 => x"e3",
  3564 => x"87",
  3565 => x"c1",
  3566 => x"cb",
  3567 => x"f6",
  3568 => x"ab",
  3569 => x"02",
  3570 => x"de",
  3571 => x"87",
  3572 => x"d8",
  3573 => x"66",
  3574 => x"4c",
  3575 => x"dc",
  3576 => x"66",
  3577 => x"1e",
  3578 => x"c1",
  3579 => x"8b",
  3580 => x"97",
  3581 => x"6b",
  3582 => x"49",
  3583 => x"74",
  3584 => x"0f",
  3585 => x"c4",
  3586 => x"86",
  3587 => x"6e",
  3588 => x"48",
  3589 => x"c1",
  3590 => x"80",
  3591 => x"c4",
  3592 => x"a6",
  3593 => x"58",
  3594 => x"c1",
  3595 => x"cb",
  3596 => x"f6",
  3597 => x"ab",
  3598 => x"05",
  3599 => x"ff",
  3600 => x"e5",
  3601 => x"87",
  3602 => x"6e",
  3603 => x"48",
  3604 => x"fc",
  3605 => x"8e",
  3606 => x"26",
  3607 => x"4d",
  3608 => x"26",
  3609 => x"4c",
  3610 => x"26",
  3611 => x"4b",
  3612 => x"26",
  3613 => x"4f",
  3614 => x"30",
  3615 => x"31",
  3616 => x"32",
  3617 => x"33",
  3618 => x"34",
  3619 => x"35",
  3620 => x"36",
  3621 => x"37",
  3622 => x"38",
  3623 => x"39",
  3624 => x"41",
  3625 => x"42",
  3626 => x"43",
  3627 => x"44",
  3628 => x"45",
  3629 => x"46",
  3630 => x"00",
  3631 => x"0e",
  3632 => x"5e",
  3633 => x"5b",
  3634 => x"5c",
  3635 => x"5d",
  3636 => x"0e",
  3637 => x"71",
  3638 => x"4b",
  3639 => x"ff",
  3640 => x"4d",
  3641 => x"13",
  3642 => x"4c",
  3643 => x"74",
  3644 => x"9c",
  3645 => x"02",
  3646 => x"d8",
  3647 => x"87",
  3648 => x"c1",
  3649 => x"85",
  3650 => x"d4",
  3651 => x"66",
  3652 => x"1e",
  3653 => x"74",
  3654 => x"49",
  3655 => x"d4",
  3656 => x"66",
  3657 => x"0f",
  3658 => x"c4",
  3659 => x"86",
  3660 => x"74",
  3661 => x"a8",
  3662 => x"05",
  3663 => x"c7",
  3664 => x"87",
  3665 => x"13",
  3666 => x"4c",
  3667 => x"74",
  3668 => x"9c",
  3669 => x"05",
  3670 => x"e8",
  3671 => x"87",
  3672 => x"75",
  3673 => x"48",
  3674 => x"26",
  3675 => x"4d",
  3676 => x"26",
  3677 => x"4c",
  3678 => x"26",
  3679 => x"4b",
  3680 => x"26",
  3681 => x"4f",
  3682 => x"0e",
  3683 => x"5e",
  3684 => x"5b",
  3685 => x"5c",
  3686 => x"5d",
  3687 => x"0e",
  3688 => x"e8",
  3689 => x"86",
  3690 => x"c4",
  3691 => x"a6",
  3692 => x"59",
  3693 => x"c0",
  3694 => x"e8",
  3695 => x"66",
  3696 => x"4d",
  3697 => x"c0",
  3698 => x"4c",
  3699 => x"c8",
  3700 => x"a6",
  3701 => x"48",
  3702 => x"c0",
  3703 => x"78",
  3704 => x"6e",
  3705 => x"97",
  3706 => x"bf",
  3707 => x"4b",
  3708 => x"6e",
  3709 => x"48",
  3710 => x"c1",
  3711 => x"80",
  3712 => x"c4",
  3713 => x"a6",
  3714 => x"58",
  3715 => x"73",
  3716 => x"9b",
  3717 => x"02",
  3718 => x"c6",
  3719 => x"d3",
  3720 => x"87",
  3721 => x"c8",
  3722 => x"66",
  3723 => x"02",
  3724 => x"c5",
  3725 => x"db",
  3726 => x"87",
  3727 => x"cc",
  3728 => x"a6",
  3729 => x"48",
  3730 => x"c0",
  3731 => x"78",
  3732 => x"fc",
  3733 => x"80",
  3734 => x"c0",
  3735 => x"78",
  3736 => x"73",
  3737 => x"4a",
  3738 => x"c0",
  3739 => x"e0",
  3740 => x"8a",
  3741 => x"02",
  3742 => x"c3",
  3743 => x"c6",
  3744 => x"87",
  3745 => x"c3",
  3746 => x"8a",
  3747 => x"02",
  3748 => x"c3",
  3749 => x"c0",
  3750 => x"87",
  3751 => x"c2",
  3752 => x"8a",
  3753 => x"02",
  3754 => x"c2",
  3755 => x"e8",
  3756 => x"87",
  3757 => x"c2",
  3758 => x"8a",
  3759 => x"02",
  3760 => x"c2",
  3761 => x"f4",
  3762 => x"87",
  3763 => x"c4",
  3764 => x"8a",
  3765 => x"02",
  3766 => x"c2",
  3767 => x"ee",
  3768 => x"87",
  3769 => x"c2",
  3770 => x"8a",
  3771 => x"02",
  3772 => x"c2",
  3773 => x"e8",
  3774 => x"87",
  3775 => x"c3",
  3776 => x"8a",
  3777 => x"02",
  3778 => x"c2",
  3779 => x"ea",
  3780 => x"87",
  3781 => x"d4",
  3782 => x"8a",
  3783 => x"02",
  3784 => x"c0",
  3785 => x"f6",
  3786 => x"87",
  3787 => x"d4",
  3788 => x"8a",
  3789 => x"02",
  3790 => x"c1",
  3791 => x"c0",
  3792 => x"87",
  3793 => x"ca",
  3794 => x"8a",
  3795 => x"02",
  3796 => x"c0",
  3797 => x"f2",
  3798 => x"87",
  3799 => x"c1",
  3800 => x"8a",
  3801 => x"02",
  3802 => x"c1",
  3803 => x"e1",
  3804 => x"87",
  3805 => x"c1",
  3806 => x"8a",
  3807 => x"02",
  3808 => x"df",
  3809 => x"87",
  3810 => x"c8",
  3811 => x"8a",
  3812 => x"02",
  3813 => x"c1",
  3814 => x"ce",
  3815 => x"87",
  3816 => x"c4",
  3817 => x"8a",
  3818 => x"02",
  3819 => x"c0",
  3820 => x"e3",
  3821 => x"87",
  3822 => x"c3",
  3823 => x"8a",
  3824 => x"02",
  3825 => x"c0",
  3826 => x"e5",
  3827 => x"87",
  3828 => x"c2",
  3829 => x"8a",
  3830 => x"02",
  3831 => x"c8",
  3832 => x"87",
  3833 => x"c3",
  3834 => x"8a",
  3835 => x"02",
  3836 => x"d3",
  3837 => x"87",
  3838 => x"c1",
  3839 => x"fa",
  3840 => x"87",
  3841 => x"cc",
  3842 => x"a6",
  3843 => x"48",
  3844 => x"ca",
  3845 => x"78",
  3846 => x"c2",
  3847 => x"d2",
  3848 => x"87",
  3849 => x"cc",
  3850 => x"a6",
  3851 => x"48",
  3852 => x"c2",
  3853 => x"78",
  3854 => x"c2",
  3855 => x"ca",
  3856 => x"87",
  3857 => x"cc",
  3858 => x"a6",
  3859 => x"48",
  3860 => x"d0",
  3861 => x"78",
  3862 => x"c2",
  3863 => x"c2",
  3864 => x"87",
  3865 => x"c0",
  3866 => x"f0",
  3867 => x"66",
  3868 => x"1e",
  3869 => x"c0",
  3870 => x"f0",
  3871 => x"66",
  3872 => x"1e",
  3873 => x"c4",
  3874 => x"85",
  3875 => x"75",
  3876 => x"4a",
  3877 => x"c4",
  3878 => x"8a",
  3879 => x"6a",
  3880 => x"49",
  3881 => x"fc",
  3882 => x"c3",
  3883 => x"87",
  3884 => x"c8",
  3885 => x"86",
  3886 => x"70",
  3887 => x"49",
  3888 => x"71",
  3889 => x"a4",
  3890 => x"4c",
  3891 => x"c1",
  3892 => x"e5",
  3893 => x"87",
  3894 => x"c8",
  3895 => x"a6",
  3896 => x"48",
  3897 => x"c1",
  3898 => x"78",
  3899 => x"c1",
  3900 => x"dd",
  3901 => x"87",
  3902 => x"c0",
  3903 => x"f0",
  3904 => x"66",
  3905 => x"1e",
  3906 => x"c4",
  3907 => x"85",
  3908 => x"75",
  3909 => x"4a",
  3910 => x"c4",
  3911 => x"8a",
  3912 => x"6a",
  3913 => x"49",
  3914 => x"c0",
  3915 => x"f0",
  3916 => x"66",
  3917 => x"0f",
  3918 => x"c4",
  3919 => x"86",
  3920 => x"c1",
  3921 => x"84",
  3922 => x"c1",
  3923 => x"c6",
  3924 => x"87",
  3925 => x"c0",
  3926 => x"f0",
  3927 => x"66",
  3928 => x"1e",
  3929 => x"c0",
  3930 => x"e5",
  3931 => x"49",
  3932 => x"c0",
  3933 => x"f0",
  3934 => x"66",
  3935 => x"0f",
  3936 => x"c4",
  3937 => x"86",
  3938 => x"c1",
  3939 => x"84",
  3940 => x"c0",
  3941 => x"f4",
  3942 => x"87",
  3943 => x"c8",
  3944 => x"a6",
  3945 => x"48",
  3946 => x"c1",
  3947 => x"78",
  3948 => x"c0",
  3949 => x"ec",
  3950 => x"87",
  3951 => x"d0",
  3952 => x"a6",
  3953 => x"48",
  3954 => x"c1",
  3955 => x"78",
  3956 => x"f8",
  3957 => x"80",
  3958 => x"c1",
  3959 => x"78",
  3960 => x"c0",
  3961 => x"e0",
  3962 => x"87",
  3963 => x"c0",
  3964 => x"f0",
  3965 => x"ab",
  3966 => x"06",
  3967 => x"da",
  3968 => x"87",
  3969 => x"c0",
  3970 => x"f9",
  3971 => x"ab",
  3972 => x"03",
  3973 => x"d4",
  3974 => x"87",
  3975 => x"d4",
  3976 => x"66",
  3977 => x"49",
  3978 => x"ca",
  3979 => x"91",
  3980 => x"73",
  3981 => x"4a",
  3982 => x"c0",
  3983 => x"f0",
  3984 => x"8a",
  3985 => x"d4",
  3986 => x"a6",
  3987 => x"48",
  3988 => x"72",
  3989 => x"a1",
  3990 => x"78",
  3991 => x"f4",
  3992 => x"80",
  3993 => x"c1",
  3994 => x"78",
  3995 => x"cc",
  3996 => x"66",
  3997 => x"02",
  3998 => x"c1",
  3999 => x"ea",
  4000 => x"87",
  4001 => x"c4",
  4002 => x"85",
  4003 => x"75",
  4004 => x"49",
  4005 => x"c4",
  4006 => x"89",
  4007 => x"a6",
  4008 => x"48",
  4009 => x"69",
  4010 => x"78",
  4011 => x"c1",
  4012 => x"e4",
  4013 => x"ab",
  4014 => x"05",
  4015 => x"d8",
  4016 => x"87",
  4017 => x"c4",
  4018 => x"66",
  4019 => x"48",
  4020 => x"c0",
  4021 => x"b7",
  4022 => x"a8",
  4023 => x"03",
  4024 => x"cf",
  4025 => x"87",
  4026 => x"c0",
  4027 => x"ed",
  4028 => x"49",
  4029 => x"f4",
  4030 => x"cf",
  4031 => x"87",
  4032 => x"c4",
  4033 => x"66",
  4034 => x"48",
  4035 => x"c0",
  4036 => x"08",
  4037 => x"88",
  4038 => x"c8",
  4039 => x"a6",
  4040 => x"58",
  4041 => x"d0",
  4042 => x"66",
  4043 => x"1e",
  4044 => x"d8",
  4045 => x"66",
  4046 => x"1e",
  4047 => x"c0",
  4048 => x"f8",
  4049 => x"66",
  4050 => x"1e",
  4051 => x"c0",
  4052 => x"f8",
  4053 => x"66",
  4054 => x"1e",
  4055 => x"dc",
  4056 => x"66",
  4057 => x"1e",
  4058 => x"d8",
  4059 => x"66",
  4060 => x"49",
  4061 => x"f6",
  4062 => x"d4",
  4063 => x"87",
  4064 => x"d4",
  4065 => x"86",
  4066 => x"70",
  4067 => x"49",
  4068 => x"71",
  4069 => x"a4",
  4070 => x"4c",
  4071 => x"c0",
  4072 => x"e1",
  4073 => x"87",
  4074 => x"c0",
  4075 => x"e5",
  4076 => x"ab",
  4077 => x"05",
  4078 => x"cf",
  4079 => x"87",
  4080 => x"d0",
  4081 => x"a6",
  4082 => x"48",
  4083 => x"c0",
  4084 => x"78",
  4085 => x"c4",
  4086 => x"80",
  4087 => x"c0",
  4088 => x"78",
  4089 => x"f4",
  4090 => x"80",
  4091 => x"c1",
  4092 => x"78",
  4093 => x"cc",
  4094 => x"87",
  4095 => x"c0",
  4096 => x"f0",
  4097 => x"66",
  4098 => x"1e",
  4099 => x"73",
  4100 => x"49",
  4101 => x"c0",
  4102 => x"f0",
  4103 => x"66",
  4104 => x"0f",
  4105 => x"c4",
  4106 => x"86",
  4107 => x"6e",
  4108 => x"97",
  4109 => x"bf",
  4110 => x"4b",
  4111 => x"6e",
  4112 => x"48",
  4113 => x"c1",
  4114 => x"80",
  4115 => x"c4",
  4116 => x"a6",
  4117 => x"58",
  4118 => x"73",
  4119 => x"9b",
  4120 => x"05",
  4121 => x"f9",
  4122 => x"ed",
  4123 => x"87",
  4124 => x"74",
  4125 => x"48",
  4126 => x"e8",
  4127 => x"8e",
  4128 => x"26",
  4129 => x"4d",
  4130 => x"26",
  4131 => x"4c",
  4132 => x"26",
  4133 => x"4b",
  4134 => x"26",
  4135 => x"4f",
  4136 => x"1e",
  4137 => x"c0",
  4138 => x"1e",
  4139 => x"c0",
  4140 => x"f3",
  4141 => x"cf",
  4142 => x"1e",
  4143 => x"d0",
  4144 => x"a6",
  4145 => x"1e",
  4146 => x"d0",
  4147 => x"66",
  4148 => x"49",
  4149 => x"f8",
  4150 => x"ea",
  4151 => x"87",
  4152 => x"f4",
  4153 => x"8e",
  4154 => x"26",
  4155 => x"4f",
  4156 => x"1e",
  4157 => x"73",
  4158 => x"1e",
  4159 => x"72",
  4160 => x"9a",
  4161 => x"02",
  4162 => x"c0",
  4163 => x"e7",
  4164 => x"87",
  4165 => x"c0",
  4166 => x"48",
  4167 => x"c1",
  4168 => x"4b",
  4169 => x"72",
  4170 => x"a9",
  4171 => x"06",
  4172 => x"d1",
  4173 => x"87",
  4174 => x"72",
  4175 => x"82",
  4176 => x"06",
  4177 => x"c9",
  4178 => x"87",
  4179 => x"73",
  4180 => x"83",
  4181 => x"72",
  4182 => x"a9",
  4183 => x"01",
  4184 => x"f4",
  4185 => x"87",
  4186 => x"c3",
  4187 => x"87",
  4188 => x"c1",
  4189 => x"b2",
  4190 => x"3a",
  4191 => x"72",
  4192 => x"a9",
  4193 => x"03",
  4194 => x"89",
  4195 => x"73",
  4196 => x"80",
  4197 => x"07",
  4198 => x"c1",
  4199 => x"2a",
  4200 => x"2b",
  4201 => x"05",
  4202 => x"f3",
  4203 => x"87",
  4204 => x"26",
  4205 => x"4b",
  4206 => x"26",
  4207 => x"4f",
  4208 => x"1e",
  4209 => x"75",
  4210 => x"1e",
  4211 => x"c4",
  4212 => x"4d",
  4213 => x"71",
  4214 => x"b7",
  4215 => x"a1",
  4216 => x"04",
  4217 => x"ff",
  4218 => x"b9",
  4219 => x"c1",
  4220 => x"81",
  4221 => x"c3",
  4222 => x"bd",
  4223 => x"07",
  4224 => x"72",
  4225 => x"b7",
  4226 => x"a2",
  4227 => x"04",
  4228 => x"ff",
  4229 => x"ba",
  4230 => x"c1",
  4231 => x"82",
  4232 => x"c1",
  4233 => x"bd",
  4234 => x"07",
  4235 => x"fe",
  4236 => x"ee",
  4237 => x"87",
  4238 => x"c1",
  4239 => x"2d",
  4240 => x"04",
  4241 => x"ff",
  4242 => x"b8",
  4243 => x"c1",
  4244 => x"80",
  4245 => x"07",
  4246 => x"2d",
  4247 => x"04",
  4248 => x"ff",
  4249 => x"b9",
  4250 => x"c1",
  4251 => x"81",
  4252 => x"07",
  4253 => x"26",
  4254 => x"4d",
  4255 => x"26",
  4256 => x"4f",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;

