library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM-2 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
type ram_type is array (0 to 2 ** (maxAddrBitBRAM-3) - 1) of word_t;

signal ram : ram_type :=
(
     0 => (x"01",x"da",x"87",x"04"),
     1 => (x"dd",x"87",x"0e",x"58"),
     2 => (x"5e",x"59",x"5a",x"0e"),
     3 => (x"27",x"00",x"00",x"00"),
     4 => (x"2c",x"0f",x"26",x"4a"),
     5 => (x"26",x"49",x"26",x"48"),
     6 => (x"ff",x"80",x"26",x"08"),
     7 => (x"4f",x"27",x"00",x"00"),
     8 => (x"00",x"2d",x"4f",x"27"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"4f",x"00",x"fd",x"87"),
    11 => (x"4f",x"c1",x"cb",x"d8"),
    12 => (x"4e",x"c9",x"c0",x"86"),
    13 => (x"c1",x"cb",x"d8",x"49"),
    14 => (x"c1",x"c1",x"f4",x"48"),
    15 => (x"89",x"d0",x"89",x"03"),
    16 => (x"c0",x"40",x"40",x"40"),
    17 => (x"40",x"f6",x"87",x"d0"),
    18 => (x"81",x"05",x"c0",x"50"),
    19 => (x"c1",x"89",x"05",x"f9"),
    20 => (x"87",x"c1",x"c1",x"f3"),
    21 => (x"4d",x"c1",x"c1",x"f3"),
    22 => (x"4c",x"74",x"ad",x"02"),
    23 => (x"c4",x"87",x"24",x"0f"),
    24 => (x"f7",x"87",x"c0",x"ec"),
    25 => (x"87",x"c1",x"c1",x"f3"),
    26 => (x"4d",x"c1",x"c1",x"f3"),
    27 => (x"4c",x"74",x"ad",x"02"),
    28 => (x"c6",x"87",x"c4",x"8c"),
    29 => (x"6c",x"0f",x"f5",x"87"),
    30 => (x"00",x"fd",x"87",x"1e"),
    31 => (x"26",x"4f",x"1e",x"73"),
    32 => (x"1e",x"c2",x"c0",x"c0"),
    33 => (x"4b",x"73",x"0f",x"c4"),
    34 => (x"87",x"26",x"4d",x"26"),
    35 => (x"4c",x"26",x"4b",x"26"),
    36 => (x"4f",x"1e",x"73",x"1e"),
    37 => (x"eb",x"48",x"c3",x"ef"),
    38 => (x"50",x"c0",x"fc",x"c0"),
    39 => (x"4b",x"c5",x"fa",x"49"),
    40 => (x"c0",x"f1",x"f9",x"87"),
    41 => (x"d1",x"c7",x"87",x"70"),
    42 => (x"98",x"02",x"c1",x"cb"),
    43 => (x"87",x"c0",x"ff",x"f0"),
    44 => (x"4b",x"c5",x"e3",x"49"),
    45 => (x"c0",x"f1",x"e5",x"87"),
    46 => (x"d6",x"fa",x"87",x"70"),
    47 => (x"98",x"02",x"c0",x"e7"),
    48 => (x"87",x"c3",x"f0",x"4b"),
    49 => (x"c2",x"c0",x"c0",x"1e"),
    50 => (x"c4",x"ca",x"49",x"c0"),
    51 => (x"ee",x"db",x"87",x"c4"),
    52 => (x"86",x"70",x"98",x"02"),
    53 => (x"c9",x"87",x"c3",x"ff"),
    54 => (x"4b",x"fe",x"e2",x"87"),
    55 => (x"c0",x"e0",x"87",x"c4"),
    56 => (x"d6",x"49",x"c0",x"f0"),
    57 => (x"f7",x"87",x"d7",x"87"),
    58 => (x"c4",x"eb",x"49",x"c0"),
    59 => (x"f0",x"ee",x"87",x"c5"),
    60 => (x"c7",x"49",x"c0",x"f0"),
    61 => (x"e7",x"87",x"c7",x"87"),
    62 => (x"c6",x"d0",x"49",x"c0"),
    63 => (x"f0",x"de",x"87",x"73"),
    64 => (x"49",x"fd",x"f7",x"87"),
    65 => (x"fe",x"d2",x"87",x"fe"),
    66 => (x"c3",x"87",x"38",x"33"),
    67 => (x"32",x"4f",x"53",x"44"),
    68 => (x"41",x"42",x"42",x"49"),
    69 => (x"4e",x"00",x"43",x"61"),
    70 => (x"6e",x"27",x"74",x"20"),
    71 => (x"6c",x"6f",x"61",x"64"),
    72 => (x"20",x"66",x"69",x"72"),
    73 => (x"6d",x"77",x"61",x"72"),
    74 => (x"65",x"0a",x"00",x"55"),
    75 => (x"6e",x"61",x"62",x"6c"),
    76 => (x"65",x"20",x"74",x"6f"),
    77 => (x"20",x"6c",x"6f",x"63"),
    78 => (x"61",x"74",x"65",x"20"),
    79 => (x"70",x"61",x"72",x"74"),
    80 => (x"69",x"74",x"69",x"6f"),
    81 => (x"6e",x"0a",x"00",x"55"),
    82 => (x"6e",x"61",x"62",x"6c"),
    83 => (x"65",x"20",x"74",x"6f"),
    84 => (x"20",x"6c",x"6f",x"63"),
    85 => (x"61",x"74",x"65",x"20"),
    86 => (x"70",x"61",x"72",x"74"),
    87 => (x"69",x"74",x"69",x"6f"),
    88 => (x"6e",x"0a",x"00",x"48"),
    89 => (x"75",x"6e",x"74",x"69"),
    90 => (x"6e",x"67",x"20",x"66"),
    91 => (x"6f",x"72",x"20",x"70"),
    92 => (x"61",x"72",x"74",x"69"),
    93 => (x"74",x"69",x"6f",x"6e"),
    94 => (x"0a",x"00",x"49",x"6e"),
    95 => (x"69",x"74",x"69",x"61"),
    96 => (x"6c",x"69",x"7a",x"69"),
    97 => (x"6e",x"67",x"20",x"53"),
    98 => (x"44",x"20",x"63",x"61"),
    99 => (x"72",x"64",x"0a",x"00"),
   100 => (x"46",x"61",x"69",x"6c"),
   101 => (x"65",x"64",x"20",x"74"),
   102 => (x"6f",x"20",x"69",x"6e"),
   103 => (x"69",x"74",x"69",x"61"),
   104 => (x"6c",x"69",x"7a",x"65"),
   105 => (x"20",x"53",x"44",x"20"),
   106 => (x"63",x"61",x"72",x"64"),
   107 => (x"0a",x"00",x"1e",x"e4"),
   108 => (x"86",x"e3",x"48",x"c3"),
   109 => (x"ff",x"50",x"e3",x"97"),
   110 => (x"bf",x"48",x"c4",x"a6"),
   111 => (x"58",x"6e",x"49",x"c3"),
   112 => (x"ff",x"99",x"e3",x"48"),
   113 => (x"c3",x"ff",x"50",x"c8"),
   114 => (x"31",x"e3",x"97",x"bf"),
   115 => (x"48",x"c8",x"a6",x"58"),
   116 => (x"c4",x"66",x"48",x"c3"),
   117 => (x"ff",x"98",x"cc",x"a6"),
   118 => (x"58",x"c8",x"66",x"b1"),
   119 => (x"e3",x"48",x"c3",x"ff"),
   120 => (x"50",x"c8",x"31",x"e3"),
   121 => (x"97",x"bf",x"48",x"d0"),
   122 => (x"a6",x"58",x"cc",x"66"),
   123 => (x"48",x"c3",x"ff",x"98"),
   124 => (x"d4",x"a6",x"58",x"d0"),
   125 => (x"66",x"b1",x"e3",x"48"),
   126 => (x"c3",x"ff",x"50",x"c8"),
   127 => (x"31",x"e3",x"97",x"bf"),
   128 => (x"48",x"d8",x"a6",x"58"),
   129 => (x"d4",x"66",x"48",x"c3"),
   130 => (x"ff",x"98",x"dc",x"a6"),
   131 => (x"58",x"d8",x"66",x"b1"),
   132 => (x"71",x"48",x"e4",x"8e"),
   133 => (x"26",x"4f",x"0e",x"5e"),
   134 => (x"5b",x"5c",x"0e",x"1e"),
   135 => (x"71",x"4a",x"72",x"49"),
   136 => (x"c3",x"ff",x"99",x"e3"),
   137 => (x"09",x"97",x"79",x"09"),
   138 => (x"c1",x"c1",x"f4",x"bf"),
   139 => (x"05",x"c8",x"87",x"d0"),
   140 => (x"66",x"48",x"c9",x"30"),
   141 => (x"d4",x"a6",x"58",x"d0"),
   142 => (x"66",x"49",x"d8",x"29"),
   143 => (x"c3",x"ff",x"99",x"e3"),
   144 => (x"09",x"97",x"79",x"09"),
   145 => (x"d0",x"66",x"49",x"d0"),
   146 => (x"29",x"c3",x"ff",x"99"),
   147 => (x"e3",x"09",x"97",x"79"),
   148 => (x"09",x"d0",x"66",x"49"),
   149 => (x"c8",x"29",x"c3",x"ff"),
   150 => (x"99",x"e3",x"09",x"97"),
   151 => (x"79",x"09",x"d0",x"66"),
   152 => (x"49",x"c3",x"ff",x"99"),
   153 => (x"e3",x"09",x"97",x"79"),
   154 => (x"09",x"72",x"49",x"d0"),
   155 => (x"29",x"c3",x"ff",x"99"),
   156 => (x"e3",x"09",x"97",x"79"),
   157 => (x"09",x"97",x"bf",x"48"),
   158 => (x"c4",x"a6",x"58",x"6e"),
   159 => (x"4b",x"c3",x"ff",x"9b"),
   160 => (x"c9",x"f0",x"ff",x"4c"),
   161 => (x"c3",x"ff",x"ab",x"05"),
   162 => (x"dc",x"87",x"e3",x"48"),
   163 => (x"c3",x"ff",x"50",x"e3"),
   164 => (x"97",x"bf",x"48",x"c4"),
   165 => (x"a6",x"58",x"6e",x"4b"),
   166 => (x"c3",x"ff",x"9b",x"c1"),
   167 => (x"8c",x"02",x"c6",x"87"),
   168 => (x"c3",x"ff",x"ab",x"02"),
   169 => (x"e4",x"87",x"73",x"4a"),
   170 => (x"c4",x"b7",x"2a",x"c0"),
   171 => (x"f0",x"a2",x"49",x"c0"),
   172 => (x"e9",x"e0",x"87",x"73"),
   173 => (x"4a",x"cf",x"9a",x"c0"),
   174 => (x"f0",x"a2",x"49",x"c0"),
   175 => (x"e9",x"d4",x"87",x"73"),
   176 => (x"48",x"26",x"c2",x"87"),
   177 => (x"26",x"4d",x"26",x"4c"),
   178 => (x"26",x"4b",x"26",x"4f"),
   179 => (x"1e",x"c0",x"49",x"e3"),
   180 => (x"48",x"c3",x"ff",x"50"),
   181 => (x"c1",x"81",x"c3",x"c8"),
   182 => (x"b7",x"a9",x"04",x"f2"),
   183 => (x"87",x"26",x"4f",x"1e"),
   184 => (x"73",x"1e",x"e8",x"87"),
   185 => (x"c4",x"f8",x"df",x"4b"),
   186 => (x"c0",x"1e",x"c0",x"ff"),
   187 => (x"f0",x"c1",x"f7",x"49"),
   188 => (x"fc",x"e3",x"87",x"c4"),
   189 => (x"86",x"c1",x"a8",x"05"),
   190 => (x"c0",x"e8",x"87",x"e3"),
   191 => (x"48",x"c3",x"ff",x"50"),
   192 => (x"c1",x"c0",x"c0",x"c0"),
   193 => (x"c0",x"c0",x"1e",x"c0"),
   194 => (x"e1",x"f0",x"c1",x"e9"),
   195 => (x"49",x"fc",x"c6",x"87"),
   196 => (x"c4",x"86",x"70",x"98"),
   197 => (x"05",x"c9",x"87",x"e3"),
   198 => (x"48",x"c3",x"ff",x"50"),
   199 => (x"c1",x"48",x"cb",x"87"),
   200 => (x"fe",x"e9",x"87",x"c1"),
   201 => (x"8b",x"05",x"fe",x"ff"),
   202 => (x"87",x"c0",x"48",x"fe"),
   203 => (x"da",x"87",x"43",x"4d"),
   204 => (x"44",x"34",x"31",x"20"),
   205 => (x"25",x"64",x"0a",x"00"),
   206 => (x"43",x"4d",x"44",x"35"),
   207 => (x"35",x"20",x"25",x"64"),
   208 => (x"0a",x"00",x"43",x"4d"),
   209 => (x"44",x"34",x"31",x"20"),
   210 => (x"25",x"64",x"0a",x"00"),
   211 => (x"43",x"4d",x"44",x"35"),
   212 => (x"35",x"20",x"25",x"64"),
   213 => (x"0a",x"00",x"69",x"6e"),
   214 => (x"69",x"74",x"20",x"25"),
   215 => (x"64",x"0a",x"20",x"20"),
   216 => (x"00",x"69",x"6e",x"69"),
   217 => (x"74",x"20",x"25",x"64"),
   218 => (x"0a",x"20",x"20",x"00"),
   219 => (x"43",x"6d",x"64",x"5f"),
   220 => (x"69",x"6e",x"69",x"74"),
   221 => (x"0a",x"00",x"43",x"4d"),
   222 => (x"44",x"38",x"5f",x"34"),
   223 => (x"20",x"72",x"65",x"73"),
   224 => (x"70",x"6f",x"6e",x"73"),
   225 => (x"65",x"3a",x"20",x"25"),
   226 => (x"64",x"0a",x"00",x"43"),
   227 => (x"4d",x"44",x"35",x"38"),
   228 => (x"20",x"25",x"64",x"0a"),
   229 => (x"20",x"20",x"00",x"43"),
   230 => (x"4d",x"44",x"35",x"38"),
   231 => (x"5f",x"32",x"20",x"25"),
   232 => (x"64",x"0a",x"20",x"20"),
   233 => (x"00",x"43",x"4d",x"44"),
   234 => (x"35",x"38",x"20",x"25"),
   235 => (x"64",x"0a",x"20",x"20"),
   236 => (x"00",x"53",x"44",x"48"),
   237 => (x"43",x"20",x"49",x"6e"),
   238 => (x"69",x"74",x"69",x"61"),
   239 => (x"6c",x"69",x"7a",x"61"),
   240 => (x"74",x"69",x"6f",x"6e"),
   241 => (x"20",x"65",x"72",x"72"),
   242 => (x"6f",x"72",x"21",x"0a"),
   243 => (x"00",x"63",x"6d",x"64"),
   244 => (x"5f",x"43",x"4d",x"44"),
   245 => (x"38",x"20",x"72",x"65"),
   246 => (x"73",x"70",x"6f",x"6e"),
   247 => (x"73",x"65",x"3a",x"20"),
   248 => (x"25",x"64",x"0a",x"00"),
   249 => (x"52",x"65",x"61",x"64"),
   250 => (x"20",x"63",x"6f",x"6d"),
   251 => (x"6d",x"61",x"6e",x"64"),
   252 => (x"20",x"66",x"61",x"69"),
   253 => (x"6c",x"65",x"64",x"20"),
   254 => (x"61",x"74",x"20",x"25"),
   255 => (x"64",x"20",x"28",x"25"),
   256 => (x"64",x"29",x"0a",x"00"),
   257 => (x"1e",x"73",x"1e",x"e3"),
   258 => (x"48",x"c3",x"ff",x"50"),
   259 => (x"cd",x"ec",x"49",x"c0"),
   260 => (x"e4",x"ca",x"87",x"d3"),
   261 => (x"4b",x"c0",x"1e",x"c0"),
   262 => (x"ff",x"f0",x"c1",x"c1"),
   263 => (x"49",x"f7",x"f6",x"87"),
   264 => (x"c4",x"86",x"70",x"98"),
   265 => (x"05",x"c9",x"87",x"e3"),
   266 => (x"48",x"c3",x"ff",x"50"),
   267 => (x"c1",x"48",x"cb",x"87"),
   268 => (x"fa",x"d9",x"87",x"c1"),
   269 => (x"8b",x"05",x"ff",x"dc"),
   270 => (x"87",x"c0",x"48",x"fa"),
   271 => (x"ca",x"87",x"1e",x"73"),
   272 => (x"1e",x"1e",x"fa",x"c7"),
   273 => (x"87",x"c6",x"ea",x"1e"),
   274 => (x"c0",x"e1",x"f0",x"c1"),
   275 => (x"c8",x"49",x"f7",x"c5"),
   276 => (x"87",x"70",x"4b",x"73"),
   277 => (x"1e",x"cf",x"cd",x"49"),
   278 => (x"c0",x"ee",x"de",x"87"),
   279 => (x"c8",x"86",x"c1",x"ab"),
   280 => (x"02",x"c8",x"87",x"fe"),
   281 => (x"de",x"87",x"c0",x"48"),
   282 => (x"c1",x"ff",x"87",x"f5"),
   283 => (x"c0",x"87",x"70",x"49"),
   284 => (x"cf",x"ff",x"ff",x"99"),
   285 => (x"c6",x"ea",x"a9",x"02"),
   286 => (x"c8",x"87",x"fe",x"c7"),
   287 => (x"87",x"c0",x"48",x"c1"),
   288 => (x"e8",x"87",x"e3",x"48"),
   289 => (x"c3",x"ff",x"50",x"c0"),
   290 => (x"f1",x"4b",x"f9",x"d2"),
   291 => (x"87",x"70",x"98",x"02"),
   292 => (x"c1",x"c6",x"87",x"c0"),
   293 => (x"1e",x"c0",x"ff",x"f0"),
   294 => (x"c1",x"fa",x"49",x"f5"),
   295 => (x"f8",x"87",x"c4",x"86"),
   296 => (x"70",x"98",x"05",x"c0"),
   297 => (x"f3",x"87",x"e3",x"48"),
   298 => (x"c3",x"ff",x"50",x"e3"),
   299 => (x"97",x"bf",x"48",x"c4"),
   300 => (x"a6",x"58",x"6e",x"49"),
   301 => (x"c3",x"ff",x"99",x"e3"),
   302 => (x"48",x"c3",x"ff",x"50"),
   303 => (x"e3",x"48",x"c3",x"ff"),
   304 => (x"50",x"e3",x"48",x"c3"),
   305 => (x"ff",x"50",x"e3",x"48"),
   306 => (x"c3",x"ff",x"50",x"c1"),
   307 => (x"c0",x"99",x"02",x"c4"),
   308 => (x"87",x"c1",x"48",x"d5"),
   309 => (x"87",x"c0",x"48",x"d1"),
   310 => (x"87",x"c2",x"ab",x"05"),
   311 => (x"c4",x"87",x"c0",x"48"),
   312 => (x"c8",x"87",x"c1",x"8b"),
   313 => (x"05",x"fe",x"e2",x"87"),
   314 => (x"c0",x"48",x"26",x"f7"),
   315 => (x"da",x"87",x"1e",x"73"),
   316 => (x"1e",x"c1",x"c1",x"f4"),
   317 => (x"48",x"c1",x"78",x"eb"),
   318 => (x"48",x"c3",x"ef",x"50"),
   319 => (x"c7",x"4b",x"e7",x"48"),
   320 => (x"c3",x"50",x"f7",x"c7"),
   321 => (x"87",x"e7",x"48",x"c2"),
   322 => (x"50",x"e3",x"48",x"c3"),
   323 => (x"ff",x"50",x"c0",x"1e"),
   324 => (x"c0",x"e5",x"d0",x"c1"),
   325 => (x"c0",x"49",x"f3",x"fd"),
   326 => (x"87",x"c4",x"86",x"c1"),
   327 => (x"a8",x"05",x"c2",x"87"),
   328 => (x"c1",x"4b",x"c2",x"ab"),
   329 => (x"05",x"c5",x"87",x"c0"),
   330 => (x"48",x"c0",x"f1",x"87"),
   331 => (x"c1",x"8b",x"05",x"ff"),
   332 => (x"cc",x"87",x"fc",x"c9"),
   333 => (x"87",x"c1",x"c1",x"f8"),
   334 => (x"58",x"c1",x"c1",x"f4"),
   335 => (x"bf",x"05",x"cd",x"87"),
   336 => (x"c1",x"1e",x"c0",x"ff"),
   337 => (x"f0",x"c1",x"d0",x"49"),
   338 => (x"f3",x"cb",x"87",x"c4"),
   339 => (x"86",x"e3",x"48",x"c3"),
   340 => (x"ff",x"50",x"e7",x"48"),
   341 => (x"c3",x"50",x"e3",x"48"),
   342 => (x"c3",x"ff",x"50",x"c1"),
   343 => (x"48",x"f5",x"e8",x"87"),
   344 => (x"0e",x"5e",x"5b",x"5c"),
   345 => (x"5d",x"0e",x"1e",x"71"),
   346 => (x"4a",x"c0",x"4d",x"e3"),
   347 => (x"48",x"c3",x"ff",x"50"),
   348 => (x"e7",x"48",x"c2",x"50"),
   349 => (x"eb",x"48",x"c7",x"50"),
   350 => (x"e3",x"48",x"c3",x"ff"),
   351 => (x"50",x"72",x"1e",x"c0"),
   352 => (x"ff",x"f0",x"c1",x"d1"),
   353 => (x"49",x"f2",x"ce",x"87"),
   354 => (x"c4",x"86",x"70",x"98"),
   355 => (x"05",x"c1",x"c9",x"87"),
   356 => (x"c5",x"ee",x"cd",x"df"),
   357 => (x"4b",x"e3",x"48",x"c3"),
   358 => (x"ff",x"50",x"e3",x"97"),
   359 => (x"bf",x"48",x"c4",x"a6"),
   360 => (x"58",x"6e",x"49",x"c3"),
   361 => (x"ff",x"99",x"c3",x"fe"),
   362 => (x"a9",x"05",x"de",x"87"),
   363 => (x"c0",x"4c",x"ef",x"fd"),
   364 => (x"87",x"d4",x"66",x"08"),
   365 => (x"78",x"08",x"d4",x"66"),
   366 => (x"48",x"c4",x"80",x"d8"),
   367 => (x"a6",x"58",x"c1",x"84"),
   368 => (x"c2",x"c0",x"b7",x"ac"),
   369 => (x"04",x"e7",x"87",x"c1"),
   370 => (x"4b",x"4d",x"c1",x"8b"),
   371 => (x"05",x"ff",x"c5",x"87"),
   372 => (x"e3",x"48",x"c3",x"ff"),
   373 => (x"50",x"e7",x"48",x"c3"),
   374 => (x"50",x"75",x"48",x"26"),
   375 => (x"f3",x"e5",x"87",x"1e"),
   376 => (x"73",x"1e",x"71",x"4b"),
   377 => (x"73",x"49",x"d8",x"29"),
   378 => (x"c3",x"ff",x"99",x"73"),
   379 => (x"4a",x"c8",x"2a",x"cf"),
   380 => (x"fc",x"c0",x"9a",x"72"),
   381 => (x"b1",x"73",x"4a",x"c8"),
   382 => (x"32",x"c0",x"ff",x"f0"),
   383 => (x"c0",x"c0",x"9a",x"72"),
   384 => (x"b1",x"73",x"4a",x"d8"),
   385 => (x"32",x"ff",x"c0",x"c0"),
   386 => (x"c0",x"c0",x"9a",x"72"),
   387 => (x"b1",x"71",x"48",x"c4"),
   388 => (x"87",x"26",x"4d",x"26"),
   389 => (x"4c",x"26",x"4b",x"26"),
   390 => (x"4f",x"1e",x"73",x"1e"),
   391 => (x"71",x"4b",x"73",x"49"),
   392 => (x"c8",x"29",x"c3",x"ff"),
   393 => (x"99",x"73",x"4a",x"c8"),
   394 => (x"32",x"cf",x"fc",x"c0"),
   395 => (x"9a",x"72",x"b1",x"71"),
   396 => (x"48",x"e2",x"87",x"0e"),
   397 => (x"5e",x"5b",x"5c",x"0e"),
   398 => (x"71",x"4b",x"c0",x"4c"),
   399 => (x"d0",x"66",x"48",x"c0"),
   400 => (x"b7",x"a8",x"06",x"c0"),
   401 => (x"e3",x"87",x"13",x"4a"),
   402 => (x"cc",x"66",x"97",x"bf"),
   403 => (x"49",x"cc",x"66",x"48"),
   404 => (x"c1",x"80",x"d0",x"a6"),
   405 => (x"58",x"71",x"b7",x"aa"),
   406 => (x"02",x"c4",x"87",x"c1"),
   407 => (x"48",x"cc",x"87",x"c1"),
   408 => (x"84",x"d0",x"66",x"b7"),
   409 => (x"ac",x"04",x"ff",x"dd"),
   410 => (x"87",x"c0",x"48",x"c2"),
   411 => (x"87",x"26",x"4d",x"26"),
   412 => (x"4c",x"26",x"4b",x"26"),
   413 => (x"4f",x"0e",x"5e",x"5b"),
   414 => (x"5c",x"0e",x"1e",x"c1"),
   415 => (x"ca",x"f6",x"48",x"ff"),
   416 => (x"78",x"c1",x"ca",x"c6"),
   417 => (x"48",x"c0",x"78",x"c0"),
   418 => (x"e7",x"da",x"49",x"da"),
   419 => (x"cf",x"87",x"c1",x"c1"),
   420 => (x"fe",x"1e",x"c0",x"49"),
   421 => (x"fb",x"c9",x"87",x"c4"),
   422 => (x"86",x"70",x"98",x"05"),
   423 => (x"c5",x"87",x"c0",x"48"),
   424 => (x"ca",x"f0",x"87",x"c0"),
   425 => (x"4b",x"c1",x"ca",x"f2"),
   426 => (x"48",x"c1",x"78",x"c8"),
   427 => (x"1e",x"c0",x"e7",x"e7"),
   428 => (x"1e",x"c1",x"c2",x"f4"),
   429 => (x"49",x"fd",x"fb",x"87"),
   430 => (x"c8",x"86",x"70",x"98"),
   431 => (x"05",x"c6",x"87",x"c1"),
   432 => (x"ca",x"f2",x"48",x"c0"),
   433 => (x"78",x"c8",x"1e",x"c0"),
   434 => (x"e7",x"f0",x"1e",x"c1"),
   435 => (x"c3",x"d0",x"49",x"fd"),
   436 => (x"e1",x"87",x"c8",x"86"),
   437 => (x"70",x"98",x"05",x"c6"),
   438 => (x"87",x"c1",x"ca",x"f2"),
   439 => (x"48",x"c0",x"78",x"c8"),
   440 => (x"1e",x"c0",x"e7",x"f9"),
   441 => (x"1e",x"c1",x"c3",x"d0"),
   442 => (x"49",x"fd",x"c7",x"87"),
   443 => (x"c8",x"86",x"70",x"98"),
   444 => (x"05",x"c5",x"87",x"c0"),
   445 => (x"48",x"c9",x"db",x"87"),
   446 => (x"c1",x"ca",x"f2",x"bf"),
   447 => (x"1e",x"c0",x"e8",x"c2"),
   448 => (x"1e",x"c0",x"e3",x"f5"),
   449 => (x"87",x"c8",x"86",x"c1"),
   450 => (x"ca",x"f2",x"bf",x"02"),
   451 => (x"c1",x"ed",x"87",x"c1"),
   452 => (x"c1",x"fe",x"4a",x"48"),
   453 => (x"c6",x"fe",x"a0",x"4c"),
   454 => (x"c1",x"c9",x"c4",x"bf"),
   455 => (x"4b",x"c1",x"c9",x"fc"),
   456 => (x"9f",x"bf",x"49",x"c4"),
   457 => (x"a6",x"5a",x"c5",x"d6"),
   458 => (x"ea",x"a9",x"05",x"c0"),
   459 => (x"cc",x"87",x"c8",x"a4"),
   460 => (x"4a",x"6a",x"49",x"fa"),
   461 => (x"e9",x"87",x"70",x"4b"),
   462 => (x"db",x"87",x"c7",x"fe"),
   463 => (x"a2",x"49",x"9f",x"69"),
   464 => (x"49",x"ca",x"e9",x"d5"),
   465 => (x"a9",x"02",x"c0",x"cc"),
   466 => (x"87",x"c0",x"e5",x"d7"),
   467 => (x"49",x"d7",x"cd",x"87"),
   468 => (x"c0",x"48",x"c7",x"fe"),
   469 => (x"87",x"73",x"1e",x"c0"),
   470 => (x"e5",x"f5",x"1e",x"c0"),
   471 => (x"e2",x"db",x"87",x"c1"),
   472 => (x"c1",x"fe",x"1e",x"73"),
   473 => (x"49",x"f7",x"f8",x"87"),
   474 => (x"cc",x"86",x"70",x"98"),
   475 => (x"05",x"c0",x"c5",x"87"),
   476 => (x"c0",x"48",x"c7",x"de"),
   477 => (x"87",x"c0",x"e6",x"cd"),
   478 => (x"49",x"d6",x"e1",x"87"),
   479 => (x"c0",x"e8",x"d5",x"1e"),
   480 => (x"c0",x"e1",x"f6",x"87"),
   481 => (x"c8",x"1e",x"c0",x"e8"),
   482 => (x"ed",x"1e",x"c1",x"c3"),
   483 => (x"d0",x"49",x"fa",x"e2"),
   484 => (x"87",x"cc",x"86",x"70"),
   485 => (x"98",x"05",x"c0",x"c9"),
   486 => (x"87",x"c1",x"ca",x"c6"),
   487 => (x"48",x"c1",x"78",x"c0"),
   488 => (x"e4",x"87",x"c8",x"1e"),
   489 => (x"c0",x"e8",x"f6",x"1e"),
   490 => (x"c1",x"c2",x"f4",x"49"),
   491 => (x"fa",x"c4",x"87",x"c8"),
   492 => (x"86",x"70",x"98",x"02"),
   493 => (x"c0",x"cf",x"87",x"c0"),
   494 => (x"e6",x"f4",x"1e",x"c0"),
   495 => (x"e0",x"fb",x"87",x"c4"),
   496 => (x"86",x"c0",x"48",x"c6"),
   497 => (x"cd",x"87",x"c1",x"c9"),
   498 => (x"fc",x"97",x"bf",x"49"),
   499 => (x"c1",x"d5",x"a9",x"05"),
   500 => (x"c0",x"cd",x"87",x"c1"),
   501 => (x"c9",x"fd",x"97",x"bf"),
   502 => (x"49",x"c2",x"ea",x"a9"),
   503 => (x"02",x"c0",x"c5",x"87"),
   504 => (x"c0",x"48",x"c5",x"ee"),
   505 => (x"87",x"c1",x"c1",x"fe"),
   506 => (x"97",x"bf",x"49",x"c3"),
   507 => (x"e9",x"a9",x"02",x"c0"),
   508 => (x"d2",x"87",x"c1",x"c1"),
   509 => (x"fe",x"97",x"bf",x"49"),
   510 => (x"c3",x"eb",x"a9",x"02"),
   511 => (x"c0",x"c5",x"87",x"c0"),
   512 => (x"48",x"c5",x"cf",x"87"),
   513 => (x"c1",x"c2",x"c9",x"97"),
   514 => (x"bf",x"49",x"71",x"99"),
   515 => (x"05",x"c0",x"cc",x"87"),
   516 => (x"c1",x"c2",x"ca",x"97"),
   517 => (x"bf",x"49",x"c2",x"a9"),
   518 => (x"02",x"c0",x"c5",x"87"),
   519 => (x"c0",x"48",x"c4",x"f2"),
   520 => (x"87",x"c1",x"c2",x"cb"),
   521 => (x"97",x"bf",x"48",x"c1"),
   522 => (x"ca",x"c2",x"58",x"c1"),
   523 => (x"c9",x"fe",x"bf",x"48"),
   524 => (x"c1",x"88",x"c1",x"ca"),
   525 => (x"c6",x"58",x"c1",x"c2"),
   526 => (x"cc",x"97",x"bf",x"49"),
   527 => (x"73",x"81",x"c1",x"c2"),
   528 => (x"cd",x"97",x"bf",x"4a"),
   529 => (x"c8",x"32",x"c1",x"ca"),
   530 => (x"d2",x"48",x"72",x"a1"),
   531 => (x"78",x"c1",x"c2",x"ce"),
   532 => (x"97",x"bf",x"48",x"c1"),
   533 => (x"ca",x"ea",x"58",x"c1"),
   534 => (x"ca",x"c6",x"bf",x"02"),
   535 => (x"c2",x"e2",x"87",x"c8"),
   536 => (x"1e",x"c0",x"e7",x"d1"),
   537 => (x"1e",x"c1",x"c3",x"d0"),
   538 => (x"49",x"f7",x"c7",x"87"),
   539 => (x"c8",x"86",x"70",x"98"),
   540 => (x"02",x"c0",x"c5",x"87"),
   541 => (x"c0",x"48",x"c3",x"da"),
   542 => (x"87",x"c1",x"c9",x"fe"),
   543 => (x"bf",x"48",x"c4",x"30"),
   544 => (x"c1",x"ca",x"ee",x"58"),
   545 => (x"c1",x"c9",x"fe",x"bf"),
   546 => (x"4a",x"c1",x"ca",x"e6"),
   547 => (x"5a",x"c1",x"c2",x"e3"),
   548 => (x"97",x"bf",x"49",x"c8"),
   549 => (x"31",x"c1",x"c2",x"e2"),
   550 => (x"97",x"bf",x"4b",x"73"),
   551 => (x"a1",x"49",x"c1",x"c2"),
   552 => (x"e4",x"97",x"bf",x"4b"),
   553 => (x"d0",x"33",x"73",x"a1"),
   554 => (x"49",x"c1",x"c2",x"e5"),
   555 => (x"97",x"bf",x"4b",x"d8"),
   556 => (x"33",x"73",x"a1",x"49"),
   557 => (x"c1",x"ca",x"f2",x"59"),
   558 => (x"c1",x"ca",x"e6",x"bf"),
   559 => (x"91",x"c1",x"ca",x"d2"),
   560 => (x"bf",x"81",x"c1",x"ca"),
   561 => (x"da",x"59",x"c1",x"c2"),
   562 => (x"eb",x"97",x"bf",x"4b"),
   563 => (x"c8",x"33",x"c1",x"c2"),
   564 => (x"ea",x"97",x"bf",x"4c"),
   565 => (x"74",x"a3",x"4b",x"c1"),
   566 => (x"c2",x"ec",x"97",x"bf"),
   567 => (x"4c",x"d0",x"34",x"74"),
   568 => (x"a3",x"4b",x"c1",x"c2"),
   569 => (x"ed",x"97",x"bf",x"4c"),
   570 => (x"cf",x"9c",x"d8",x"34"),
   571 => (x"74",x"a3",x"4b",x"c1"),
   572 => (x"ca",x"de",x"5b",x"c2"),
   573 => (x"8b",x"73",x"92",x"c1"),
   574 => (x"ca",x"de",x"48",x"72"),
   575 => (x"a1",x"78",x"c1",x"d0"),
   576 => (x"87",x"c1",x"c2",x"d0"),
   577 => (x"97",x"bf",x"49",x"c8"),
   578 => (x"31",x"c1",x"c2",x"cf"),
   579 => (x"97",x"bf",x"4a",x"72"),
   580 => (x"a1",x"49",x"c1",x"ca"),
   581 => (x"ee",x"59",x"c5",x"31"),
   582 => (x"c7",x"ff",x"81",x"c9"),
   583 => (x"29",x"c1",x"ca",x"e6"),
   584 => (x"59",x"c1",x"c2",x"d5"),
   585 => (x"97",x"bf",x"4a",x"c8"),
   586 => (x"32",x"c1",x"c2",x"d4"),
   587 => (x"97",x"bf",x"4b",x"73"),
   588 => (x"a2",x"4a",x"c1",x"ca"),
   589 => (x"f2",x"5a",x"c1",x"ca"),
   590 => (x"e6",x"bf",x"92",x"c1"),
   591 => (x"ca",x"d2",x"bf",x"82"),
   592 => (x"c1",x"ca",x"e2",x"5a"),
   593 => (x"c1",x"ca",x"da",x"48"),
   594 => (x"c0",x"78",x"c1",x"ca"),
   595 => (x"d6",x"48",x"72",x"a1"),
   596 => (x"78",x"c1",x"48",x"26"),
   597 => (x"f4",x"d8",x"87",x"4e"),
   598 => (x"6f",x"20",x"70",x"61"),
   599 => (x"72",x"74",x"69",x"74"),
   600 => (x"69",x"6f",x"6e",x"20"),
   601 => (x"73",x"69",x"67",x"6e"),
   602 => (x"61",x"74",x"75",x"72"),
   603 => (x"65",x"20",x"66",x"6f"),
   604 => (x"75",x"6e",x"64",x"0a"),
   605 => (x"00",x"52",x"65",x"61"),
   606 => (x"64",x"69",x"6e",x"67"),
   607 => (x"20",x"62",x"6f",x"6f"),
   608 => (x"74",x"20",x"73",x"65"),
   609 => (x"63",x"74",x"6f",x"72"),
   610 => (x"20",x"25",x"64",x"0a"),
   611 => (x"00",x"52",x"65",x"61"),
   612 => (x"64",x"20",x"62",x"6f"),
   613 => (x"6f",x"74",x"20",x"73"),
   614 => (x"65",x"63",x"74",x"6f"),
   615 => (x"72",x"20",x"66",x"72"),
   616 => (x"6f",x"6d",x"20",x"66"),
   617 => (x"69",x"72",x"73",x"74"),
   618 => (x"20",x"70",x"61",x"72"),
   619 => (x"74",x"69",x"74",x"69"),
   620 => (x"6f",x"6e",x"0a",x"00"),
   621 => (x"55",x"6e",x"73",x"75"),
   622 => (x"70",x"70",x"6f",x"72"),
   623 => (x"74",x"65",x"64",x"20"),
   624 => (x"70",x"61",x"72",x"74"),
   625 => (x"69",x"74",x"69",x"6f"),
   626 => (x"6e",x"20",x"74",x"79"),
   627 => (x"70",x"65",x"21",x"0d"),
   628 => (x"00",x"46",x"41",x"54"),
   629 => (x"33",x"32",x"20",x"20"),
   630 => (x"20",x"00",x"52",x"65"),
   631 => (x"61",x"64",x"69",x"6e"),
   632 => (x"67",x"20",x"4d",x"42"),
   633 => (x"52",x"0a",x"00",x"46"),
   634 => (x"41",x"54",x"31",x"36"),
   635 => (x"20",x"20",x"20",x"00"),
   636 => (x"46",x"41",x"54",x"33"),
   637 => (x"32",x"20",x"20",x"20"),
   638 => (x"00",x"46",x"41",x"54"),
   639 => (x"31",x"32",x"20",x"20"),
   640 => (x"20",x"00",x"50",x"61"),
   641 => (x"72",x"74",x"69",x"74"),
   642 => (x"69",x"6f",x"6e",x"63"),
   643 => (x"6f",x"75",x"6e",x"74"),
   644 => (x"20",x"25",x"64",x"0a"),
   645 => (x"00",x"48",x"75",x"6e"),
   646 => (x"74",x"69",x"6e",x"67"),
   647 => (x"20",x"66",x"6f",x"72"),
   648 => (x"20",x"66",x"69",x"6c"),
   649 => (x"65",x"73",x"79",x"73"),
   650 => (x"74",x"65",x"6d",x"0a"),
   651 => (x"00",x"46",x"41",x"54"),
   652 => (x"33",x"32",x"20",x"20"),
   653 => (x"20",x"00",x"46",x"41"),
   654 => (x"54",x"31",x"36",x"20"),
   655 => (x"20",x"20",x"00",x"52"),
   656 => (x"65",x"61",x"64",x"69"),
   657 => (x"6e",x"67",x"20",x"64"),
   658 => (x"69",x"72",x"65",x"63"),
   659 => (x"74",x"6f",x"72",x"79"),
   660 => (x"20",x"73",x"65",x"63"),
   661 => (x"74",x"6f",x"72",x"20"),
   662 => (x"25",x"64",x"0a",x"00"),
   663 => (x"66",x"69",x"6c",x"65"),
   664 => (x"20",x"22",x"25",x"73"),
   665 => (x"22",x"20",x"66",x"6f"),
   666 => (x"75",x"6e",x"64",x"0d"),
   667 => (x"00",x"47",x"65",x"74"),
   668 => (x"46",x"41",x"54",x"4c"),
   669 => (x"69",x"6e",x"6b",x"20"),
   670 => (x"72",x"65",x"74",x"75"),
   671 => (x"72",x"6e",x"65",x"64"),
   672 => (x"20",x"25",x"64",x"0a"),
   673 => (x"00",x"43",x"61",x"6e"),
   674 => (x"27",x"74",x"20",x"6f"),
   675 => (x"70",x"65",x"6e",x"20"),
   676 => (x"25",x"73",x"0a",x"00"),
   677 => (x"0e",x"5e",x"5b",x"5c"),
   678 => (x"5d",x"0e",x"71",x"4a"),
   679 => (x"c1",x"ca",x"c6",x"bf"),
   680 => (x"02",x"cc",x"87",x"72"),
   681 => (x"4b",x"c7",x"b7",x"2b"),
   682 => (x"72",x"4c",x"c1",x"ff"),
   683 => (x"9c",x"ca",x"87",x"72"),
   684 => (x"4b",x"c8",x"b7",x"2b"),
   685 => (x"72",x"4c",x"c3",x"ff"),
   686 => (x"9c",x"c1",x"ca",x"f6"),
   687 => (x"bf",x"ab",x"02",x"de"),
   688 => (x"87",x"c1",x"c1",x"fe"),
   689 => (x"1e",x"c1",x"ca",x"d2"),
   690 => (x"bf",x"49",x"73",x"81"),
   691 => (x"ea",x"d1",x"87",x"c4"),
   692 => (x"86",x"70",x"98",x"05"),
   693 => (x"c5",x"87",x"c0",x"48"),
   694 => (x"c0",x"f6",x"87",x"c1"),
   695 => (x"ca",x"fa",x"5b",x"c1"),
   696 => (x"ca",x"c6",x"bf",x"02"),
   697 => (x"d9",x"87",x"74",x"4a"),
   698 => (x"c4",x"92",x"c1",x"c1"),
   699 => (x"fe",x"82",x"6a",x"49"),
   700 => (x"eb",x"ec",x"87",x"70"),
   701 => (x"49",x"71",x"4d",x"cf"),
   702 => (x"ff",x"ff",x"ff",x"ff"),
   703 => (x"9d",x"d0",x"87",x"74"),
   704 => (x"4a",x"c2",x"92",x"c1"),
   705 => (x"c1",x"fe",x"82",x"9f"),
   706 => (x"6a",x"49",x"ec",x"cc"),
   707 => (x"87",x"70",x"4d",x"75"),
   708 => (x"48",x"ed",x"d9",x"87"),
   709 => (x"0e",x"5e",x"5b",x"5c"),
   710 => (x"5d",x"0e",x"f4",x"86"),
   711 => (x"71",x"4c",x"c0",x"4b"),
   712 => (x"c1",x"ca",x"f6",x"48"),
   713 => (x"ff",x"78",x"c1",x"ca"),
   714 => (x"da",x"bf",x"4d",x"c1"),
   715 => (x"ca",x"de",x"bf",x"7e"),
   716 => (x"c1",x"ca",x"c6",x"bf"),
   717 => (x"02",x"c9",x"87",x"c1"),
   718 => (x"c9",x"fe",x"bf",x"4a"),
   719 => (x"c4",x"32",x"c7",x"87"),
   720 => (x"c1",x"ca",x"e2",x"bf"),
   721 => (x"4a",x"c4",x"32",x"c8"),
   722 => (x"a6",x"5a",x"c8",x"a6"),
   723 => (x"48",x"c0",x"78",x"c4"),
   724 => (x"66",x"48",x"c0",x"a8"),
   725 => (x"06",x"c3",x"cf",x"87"),
   726 => (x"c8",x"66",x"49",x"cf"),
   727 => (x"99",x"05",x"c0",x"e3"),
   728 => (x"87",x"6e",x"1e",x"c0"),
   729 => (x"e8",x"ff",x"1e",x"d2"),
   730 => (x"d0",x"87",x"c1",x"c1"),
   731 => (x"fe",x"1e",x"cc",x"66"),
   732 => (x"49",x"48",x"c1",x"80"),
   733 => (x"d0",x"a6",x"58",x"71"),
   734 => (x"49",x"e7",x"e4",x"87"),
   735 => (x"cc",x"86",x"c1",x"c1"),
   736 => (x"fe",x"4b",x"c3",x"87"),
   737 => (x"c0",x"e0",x"83",x"97"),
   738 => (x"6b",x"49",x"71",x"99"),
   739 => (x"02",x"c2",x"c5",x"87"),
   740 => (x"97",x"6b",x"49",x"c3"),
   741 => (x"e5",x"a9",x"02",x"c1"),
   742 => (x"fb",x"87",x"cb",x"a3"),
   743 => (x"49",x"97",x"69",x"49"),
   744 => (x"d8",x"99",x"05",x"c1"),
   745 => (x"ef",x"87",x"cb",x"1e"),
   746 => (x"c0",x"e0",x"66",x"1e"),
   747 => (x"73",x"49",x"ea",x"c2"),
   748 => (x"87",x"c8",x"86",x"70"),
   749 => (x"98",x"05",x"c1",x"dc"),
   750 => (x"87",x"dc",x"a3",x"4a"),
   751 => (x"6a",x"49",x"e8",x"de"),
   752 => (x"87",x"70",x"4a",x"c4"),
   753 => (x"a4",x"49",x"72",x"79"),
   754 => (x"da",x"a3",x"4a",x"9f"),
   755 => (x"6a",x"49",x"e9",x"c8"),
   756 => (x"87",x"c4",x"a6",x"58"),
   757 => (x"c1",x"ca",x"c6",x"bf"),
   758 => (x"02",x"d8",x"87",x"d4"),
   759 => (x"a3",x"4a",x"9f",x"6a"),
   760 => (x"49",x"e8",x"f5",x"87"),
   761 => (x"70",x"49",x"c0",x"ff"),
   762 => (x"ff",x"99",x"71",x"48"),
   763 => (x"d0",x"30",x"c8",x"a6"),
   764 => (x"58",x"c5",x"87",x"c4"),
   765 => (x"a6",x"48",x"c0",x"78"),
   766 => (x"c4",x"66",x"4a",x"6e"),
   767 => (x"82",x"c8",x"a4",x"49"),
   768 => (x"72",x"79",x"c0",x"7c"),
   769 => (x"dc",x"66",x"1e",x"c0"),
   770 => (x"e9",x"dc",x"1e",x"cf"),
   771 => (x"ec",x"87",x"c8",x"86"),
   772 => (x"c1",x"48",x"c1",x"d0"),
   773 => (x"87",x"c8",x"66",x"48"),
   774 => (x"c1",x"80",x"cc",x"a6"),
   775 => (x"58",x"c8",x"66",x"48"),
   776 => (x"c4",x"66",x"a8",x"04"),
   777 => (x"fc",x"f1",x"87",x"c1"),
   778 => (x"ca",x"c6",x"bf",x"02"),
   779 => (x"c0",x"f4",x"87",x"75"),
   780 => (x"49",x"f9",x"e0",x"87"),
   781 => (x"70",x"4d",x"75",x"1e"),
   782 => (x"c0",x"e9",x"ed",x"1e"),
   783 => (x"ce",x"fb",x"87",x"c8"),
   784 => (x"86",x"75",x"49",x"cf"),
   785 => (x"ff",x"ff",x"ff",x"f8"),
   786 => (x"99",x"a9",x"02",x"d6"),
   787 => (x"87",x"75",x"49",x"c2"),
   788 => (x"89",x"c1",x"c9",x"fe"),
   789 => (x"bf",x"91",x"c1",x"ca"),
   790 => (x"d6",x"bf",x"48",x"71"),
   791 => (x"80",x"c4",x"a6",x"58"),
   792 => (x"fb",x"e7",x"87",x"c0"),
   793 => (x"48",x"f4",x"8e",x"e8"),
   794 => (x"c3",x"87",x"0e",x"5e"),
   795 => (x"5b",x"5c",x"5d",x"0e"),
   796 => (x"1e",x"71",x"4b",x"73"),
   797 => (x"1e",x"c1",x"ca",x"fa"),
   798 => (x"49",x"fa",x"d8",x"87"),
   799 => (x"c4",x"86",x"70",x"98"),
   800 => (x"02",x"c1",x"f7",x"87"),
   801 => (x"c1",x"ca",x"fe",x"bf"),
   802 => (x"49",x"c7",x"ff",x"81"),
   803 => (x"c9",x"29",x"c4",x"a6"),
   804 => (x"59",x"c0",x"4d",x"4c"),
   805 => (x"6e",x"48",x"c0",x"b7"),
   806 => (x"a8",x"06",x"c1",x"ed"),
   807 => (x"87",x"c1",x"ca",x"d6"),
   808 => (x"bf",x"49",x"c1",x"cb"),
   809 => (x"c2",x"bf",x"4a",x"c2"),
   810 => (x"8a",x"c1",x"c9",x"fe"),
   811 => (x"bf",x"92",x"72",x"a1"),
   812 => (x"49",x"c1",x"ca",x"c2"),
   813 => (x"bf",x"4a",x"74",x"9a"),
   814 => (x"72",x"a1",x"49",x"d4"),
   815 => (x"66",x"1e",x"71",x"49"),
   816 => (x"e2",x"dd",x"87",x"c4"),
   817 => (x"86",x"70",x"98",x"05"),
   818 => (x"c5",x"87",x"c0",x"48"),
   819 => (x"c1",x"c0",x"87",x"c1"),
   820 => (x"84",x"c1",x"ca",x"c2"),
   821 => (x"bf",x"49",x"74",x"99"),
   822 => (x"05",x"cc",x"87",x"c1"),
   823 => (x"cb",x"c2",x"bf",x"49"),
   824 => (x"f6",x"f1",x"87",x"c1"),
   825 => (x"cb",x"c6",x"58",x"d4"),
   826 => (x"66",x"48",x"c8",x"c0"),
   827 => (x"80",x"d8",x"a6",x"58"),
   828 => (x"c1",x"85",x"6e",x"b7"),
   829 => (x"ad",x"04",x"fe",x"e4"),
   830 => (x"87",x"cf",x"87",x"73"),
   831 => (x"1e",x"c0",x"ea",x"c5"),
   832 => (x"1e",x"cb",x"f6",x"87"),
   833 => (x"c8",x"86",x"c0",x"48"),
   834 => (x"c5",x"87",x"c1",x"ca"),
   835 => (x"fe",x"bf",x"48",x"26"),
   836 => (x"e5",x"da",x"87",x"1e"),
   837 => (x"f3",x"09",x"97",x"79"),
   838 => (x"09",x"71",x"48",x"26"),
   839 => (x"4f",x"0e",x"5e",x"5b"),
   840 => (x"5c",x"0e",x"71",x"4b"),
   841 => (x"c0",x"4c",x"13",x"4a"),
   842 => (x"72",x"9a",x"02",x"cd"),
   843 => (x"87",x"72",x"49",x"e2"),
   844 => (x"87",x"c1",x"84",x"13"),
   845 => (x"4a",x"72",x"9a",x"05"),
   846 => (x"f3",x"87",x"74",x"48"),
   847 => (x"c2",x"87",x"26",x"4d"),
   848 => (x"26",x"4c",x"26",x"4b"),
   849 => (x"26",x"4f",x"0e",x"5e"),
   850 => (x"5b",x"5c",x"5d",x"0e"),
   851 => (x"fc",x"86",x"71",x"4a"),
   852 => (x"c0",x"e0",x"66",x"4c"),
   853 => (x"c1",x"cb",x"c6",x"4b"),
   854 => (x"c0",x"7e",x"72",x"9a"),
   855 => (x"05",x"ce",x"87",x"c1"),
   856 => (x"cb",x"c7",x"4b",x"c1"),
   857 => (x"cb",x"c6",x"48",x"c0"),
   858 => (x"f0",x"50",x"c1",x"d2"),
   859 => (x"87",x"72",x"9a",x"02"),
   860 => (x"c0",x"e9",x"87",x"d4"),
   861 => (x"66",x"4d",x"72",x"1e"),
   862 => (x"72",x"49",x"75",x"4a"),
   863 => (x"ca",x"cf",x"87",x"26"),
   864 => (x"4a",x"c0",x"f7",x"f0"),
   865 => (x"81",x"11",x"53",x"71"),
   866 => (x"1e",x"72",x"49",x"75"),
   867 => (x"4a",x"c9",x"fe",x"87"),
   868 => (x"70",x"4a",x"26",x"49"),
   869 => (x"c1",x"8c",x"72",x"9a"),
   870 => (x"05",x"ff",x"da",x"87"),
   871 => (x"c0",x"b7",x"ac",x"06"),
   872 => (x"dd",x"87",x"c0",x"e4"),
   873 => (x"66",x"02",x"c5",x"87"),
   874 => (x"c0",x"f0",x"4a",x"c3"),
   875 => (x"87",x"c0",x"e0",x"4a"),
   876 => (x"73",x"0a",x"97",x"7a"),
   877 => (x"0a",x"c1",x"83",x"8c"),
   878 => (x"c0",x"b7",x"ac",x"01"),
   879 => (x"ff",x"e3",x"87",x"c1"),
   880 => (x"cb",x"c6",x"ab",x"02"),
   881 => (x"de",x"87",x"d8",x"66"),
   882 => (x"4c",x"dc",x"66",x"1e"),
   883 => (x"c1",x"8b",x"97",x"6b"),
   884 => (x"49",x"74",x"0f",x"c4"),
   885 => (x"86",x"6e",x"48",x"c1"),
   886 => (x"80",x"c4",x"a6",x"58"),
   887 => (x"c1",x"cb",x"c6",x"ab"),
   888 => (x"05",x"ff",x"e5",x"87"),
   889 => (x"6e",x"48",x"fc",x"8e"),
   890 => (x"26",x"4d",x"26",x"4c"),
   891 => (x"26",x"4b",x"26",x"4f"),
   892 => (x"30",x"31",x"32",x"33"),
   893 => (x"34",x"35",x"36",x"37"),
   894 => (x"38",x"39",x"41",x"42"),
   895 => (x"43",x"44",x"45",x"46"),
   896 => (x"00",x"0e",x"5e",x"5b"),
   897 => (x"5c",x"5d",x"0e",x"71"),
   898 => (x"4b",x"ff",x"4d",x"13"),
   899 => (x"4c",x"74",x"9c",x"02"),
   900 => (x"d8",x"87",x"c1",x"85"),
   901 => (x"d4",x"66",x"1e",x"74"),
   902 => (x"49",x"d4",x"66",x"0f"),
   903 => (x"c4",x"86",x"74",x"a8"),
   904 => (x"05",x"c7",x"87",x"13"),
   905 => (x"4c",x"74",x"9c",x"05"),
   906 => (x"e8",x"87",x"75",x"48"),
   907 => (x"26",x"4d",x"26",x"4c"),
   908 => (x"26",x"4b",x"26",x"4f"),
   909 => (x"0e",x"5e",x"5b",x"5c"),
   910 => (x"5d",x"0e",x"e8",x"86"),
   911 => (x"c4",x"a6",x"59",x"c0"),
   912 => (x"e8",x"66",x"4d",x"c0"),
   913 => (x"4c",x"c8",x"a6",x"48"),
   914 => (x"c0",x"78",x"6e",x"97"),
   915 => (x"bf",x"4b",x"6e",x"48"),
   916 => (x"c1",x"80",x"c4",x"a6"),
   917 => (x"58",x"73",x"9b",x"02"),
   918 => (x"c6",x"d3",x"87",x"c8"),
   919 => (x"66",x"02",x"c5",x"db"),
   920 => (x"87",x"cc",x"a6",x"48"),
   921 => (x"c0",x"78",x"fc",x"80"),
   922 => (x"c0",x"78",x"73",x"4a"),
   923 => (x"c0",x"e0",x"8a",x"02"),
   924 => (x"c3",x"c6",x"87",x"c3"),
   925 => (x"8a",x"02",x"c3",x"c0"),
   926 => (x"87",x"c2",x"8a",x"02"),
   927 => (x"c2",x"e8",x"87",x"c2"),
   928 => (x"8a",x"02",x"c2",x"f4"),
   929 => (x"87",x"c4",x"8a",x"02"),
   930 => (x"c2",x"ee",x"87",x"c2"),
   931 => (x"8a",x"02",x"c2",x"e8"),
   932 => (x"87",x"c3",x"8a",x"02"),
   933 => (x"c2",x"ea",x"87",x"d4"),
   934 => (x"8a",x"02",x"c0",x"f6"),
   935 => (x"87",x"d4",x"8a",x"02"),
   936 => (x"c1",x"c0",x"87",x"ca"),
   937 => (x"8a",x"02",x"c0",x"f2"),
   938 => (x"87",x"c1",x"8a",x"02"),
   939 => (x"c1",x"e1",x"87",x"c1"),
   940 => (x"8a",x"02",x"df",x"87"),
   941 => (x"c8",x"8a",x"02",x"c1"),
   942 => (x"ce",x"87",x"c4",x"8a"),
   943 => (x"02",x"c0",x"e3",x"87"),
   944 => (x"c3",x"8a",x"02",x"c0"),
   945 => (x"e5",x"87",x"c2",x"8a"),
   946 => (x"02",x"c8",x"87",x"c3"),
   947 => (x"8a",x"02",x"d3",x"87"),
   948 => (x"c1",x"fa",x"87",x"cc"),
   949 => (x"a6",x"48",x"ca",x"78"),
   950 => (x"c2",x"d2",x"87",x"cc"),
   951 => (x"a6",x"48",x"c2",x"78"),
   952 => (x"c2",x"ca",x"87",x"cc"),
   953 => (x"a6",x"48",x"d0",x"78"),
   954 => (x"c2",x"c2",x"87",x"c0"),
   955 => (x"f0",x"66",x"1e",x"c0"),
   956 => (x"f0",x"66",x"1e",x"c4"),
   957 => (x"85",x"75",x"4a",x"c4"),
   958 => (x"8a",x"6a",x"49",x"fc"),
   959 => (x"c3",x"87",x"c8",x"86"),
   960 => (x"70",x"49",x"71",x"a4"),
   961 => (x"4c",x"c1",x"e5",x"87"),
   962 => (x"c8",x"a6",x"48",x"c1"),
   963 => (x"78",x"c1",x"dd",x"87"),
   964 => (x"c0",x"f0",x"66",x"1e"),
   965 => (x"c4",x"85",x"75",x"4a"),
   966 => (x"c4",x"8a",x"6a",x"49"),
   967 => (x"c0",x"f0",x"66",x"0f"),
   968 => (x"c4",x"86",x"c1",x"84"),
   969 => (x"c1",x"c6",x"87",x"c0"),
   970 => (x"f0",x"66",x"1e",x"c0"),
   971 => (x"e5",x"49",x"c0",x"f0"),
   972 => (x"66",x"0f",x"c4",x"86"),
   973 => (x"c1",x"84",x"c0",x"f4"),
   974 => (x"87",x"c8",x"a6",x"48"),
   975 => (x"c1",x"78",x"c0",x"ec"),
   976 => (x"87",x"d0",x"a6",x"48"),
   977 => (x"c1",x"78",x"f8",x"80"),
   978 => (x"c1",x"78",x"c0",x"e0"),
   979 => (x"87",x"c0",x"f0",x"ab"),
   980 => (x"06",x"da",x"87",x"c0"),
   981 => (x"f9",x"ab",x"03",x"d4"),
   982 => (x"87",x"d4",x"66",x"49"),
   983 => (x"ca",x"91",x"73",x"4a"),
   984 => (x"c0",x"f0",x"8a",x"d4"),
   985 => (x"a6",x"48",x"72",x"a1"),
   986 => (x"78",x"f4",x"80",x"c1"),
   987 => (x"78",x"cc",x"66",x"02"),
   988 => (x"c1",x"ea",x"87",x"c4"),
   989 => (x"85",x"75",x"49",x"c4"),
   990 => (x"89",x"a6",x"48",x"69"),
   991 => (x"78",x"c1",x"e4",x"ab"),
   992 => (x"05",x"d8",x"87",x"c4"),
   993 => (x"66",x"48",x"c0",x"b7"),
   994 => (x"a8",x"03",x"cf",x"87"),
   995 => (x"c0",x"ed",x"49",x"f6"),
   996 => (x"c1",x"87",x"c4",x"66"),
   997 => (x"48",x"c0",x"08",x"88"),
   998 => (x"c8",x"a6",x"58",x"d0"),
   999 => (x"66",x"1e",x"d8",x"66"),
  1000 => (x"1e",x"c0",x"f8",x"66"),
  1001 => (x"1e",x"c0",x"f8",x"66"),
  1002 => (x"1e",x"dc",x"66",x"1e"),
  1003 => (x"d8",x"66",x"49",x"f6"),
  1004 => (x"d4",x"87",x"d4",x"86"),
  1005 => (x"70",x"49",x"71",x"a4"),
  1006 => (x"4c",x"c0",x"e1",x"87"),
  1007 => (x"c0",x"e5",x"ab",x"05"),
  1008 => (x"cf",x"87",x"d0",x"a6"),
  1009 => (x"48",x"c0",x"78",x"c4"),
  1010 => (x"80",x"c0",x"78",x"f4"),
  1011 => (x"80",x"c1",x"78",x"cc"),
  1012 => (x"87",x"c0",x"f0",x"66"),
  1013 => (x"1e",x"73",x"49",x"c0"),
  1014 => (x"f0",x"66",x"0f",x"c4"),
  1015 => (x"86",x"6e",x"97",x"bf"),
  1016 => (x"4b",x"6e",x"48",x"c1"),
  1017 => (x"80",x"c4",x"a6",x"58"),
  1018 => (x"73",x"9b",x"05",x"f9"),
  1019 => (x"ed",x"87",x"74",x"48"),
  1020 => (x"e8",x"8e",x"26",x"4d"),
  1021 => (x"26",x"4c",x"26",x"4b"),
  1022 => (x"26",x"4f",x"1e",x"c0"),
  1023 => (x"1e",x"c0",x"f4",x"d3"),
  1024 => (x"1e",x"d0",x"a6",x"1e"),
  1025 => (x"d0",x"66",x"49",x"f8"),
  1026 => (x"ea",x"87",x"f4",x"8e"),
  1027 => (x"26",x"4f",x"1e",x"73"),
  1028 => (x"1e",x"72",x"9a",x"02"),
  1029 => (x"c0",x"e7",x"87",x"c0"),
  1030 => (x"48",x"c1",x"4b",x"72"),
  1031 => (x"a9",x"06",x"d1",x"87"),
  1032 => (x"72",x"82",x"06",x"c9"),
  1033 => (x"87",x"73",x"83",x"72"),
  1034 => (x"a9",x"01",x"f4",x"87"),
  1035 => (x"c3",x"87",x"c1",x"b2"),
  1036 => (x"3a",x"72",x"a9",x"03"),
  1037 => (x"89",x"73",x"80",x"07"),
  1038 => (x"c1",x"2a",x"2b",x"05"),
  1039 => (x"f3",x"87",x"26",x"4b"),
  1040 => (x"26",x"4f",x"1e",x"75"),
  1041 => (x"1e",x"c4",x"4d",x"71"),
  1042 => (x"b7",x"a1",x"04",x"ff"),
  1043 => (x"b9",x"c1",x"81",x"c3"),
  1044 => (x"bd",x"07",x"72",x"b7"),
  1045 => (x"a2",x"04",x"ff",x"ba"),
  1046 => (x"c1",x"82",x"c1",x"bd"),
  1047 => (x"07",x"fe",x"ee",x"87"),
  1048 => (x"c1",x"2d",x"04",x"ff"),
  1049 => (x"b8",x"c1",x"80",x"07"),
  1050 => (x"2d",x"04",x"ff",x"b9"),
  1051 => (x"c1",x"81",x"07",x"26"),
  1052 => (x"4d",x"26",x"4f",x"26"),
	others => (others => x"00")
);

-- Xilinx XST attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "no_rw_check";

-- Altera Quartus attributes
attribute ramstyle: string;
attribute ramstyle of ram: signal is "no_rw_check";

signal q_local : word_t;

begin
    
	process(clk,q_local)
	begin

		q(31 downto 24)<=q_local(0);
		q(23 downto 16)<=q_local(1);
		q(15 downto 8)<=q_local(2);
		q(7 downto 0)<=q_local(3);

		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel(3) = '1') then
					ram(to_integer(unsigned(addr)))(3) <= d(7 downto 0);
				end if;
				if bytesel(2) = '1' then
					ram(to_integer(unsigned(addr)))(2) <= d(15 downto 8);
				end if;
				if bytesel(1) = '1' then
					ram(to_integer(unsigned(addr)))(1) <= d(23 downto 16);
				end if;
				if bytesel(0) = '1' then
					ram(to_integer(unsigned(addr)))(0) <= d(31 downto 24);
				end if;
			end if;
			q_local <= ram(to_integer(unsigned(addr)));
		end if;
	end process;

end arch;

