library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM-2 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111";
	-- Second port
	addr2 : in std_logic_vector(maxAddrBitBRAM-2 downto 0) := (others=>'0');
	q2 : out std_logic_vector(31 downto 0);
	d2 : in std_logic_vector(31 downto 0) := X"00000000";
	we2 : in std_logic := '0';
	bytesel2 : in std_logic_vector(3 downto 0) := "1111"	
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
type ram_type is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

signal ram : ram_type :=
(
     0 => (x"01",x"da",x"87",x"04"),
     1 => (x"dd",x"87",x"0e",x"58"),
     2 => (x"5e",x"59",x"5a",x"0e"),
     3 => (x"27",x"00",x"00",x"00"),
     4 => (x"29",x"0f",x"26",x"4a"),
     5 => (x"26",x"49",x"26",x"48"),
     6 => (x"ff",x"80",x"26",x"08"),
     7 => (x"4f",x"27",x"00",x"00"),
     8 => (x"00",x"2d",x"4f",x"27"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"4f",x"4f",x"00",x"fd"),
    11 => (x"87",x"c1",x"c9",x"f8"),
    12 => (x"4e",x"c9",x"c0",x"48"),
    13 => (x"c2",x"28",x"c1",x"d5"),
    14 => (x"ea",x"e5",x"d6",x"ea"),
    15 => (x"49",x"71",x"46",x"c1"),
    16 => (x"88",x"01",x"f9",x"87"),
    17 => (x"c1",x"c9",x"f8",x"49"),
    18 => (x"c1",x"c0",x"e4",x"48"),
    19 => (x"89",x"d0",x"89",x"03"),
    20 => (x"c0",x"40",x"40",x"40"),
    21 => (x"40",x"f6",x"87",x"d0"),
    22 => (x"81",x"05",x"c0",x"50"),
    23 => (x"c1",x"89",x"05",x"f9"),
    24 => (x"87",x"c1",x"c0",x"e2"),
    25 => (x"4d",x"c1",x"c0",x"e2"),
    26 => (x"4c",x"74",x"ad",x"02"),
    27 => (x"c4",x"87",x"24",x"0f"),
    28 => (x"f7",x"87",x"c2",x"db"),
    29 => (x"87",x"c1",x"c0",x"e2"),
    30 => (x"4d",x"c1",x"c0",x"e2"),
    31 => (x"4c",x"74",x"ad",x"02"),
    32 => (x"c6",x"87",x"c4",x"8c"),
    33 => (x"6c",x"0f",x"f5",x"87"),
    34 => (x"00",x"fd",x"87",x"0e"),
    35 => (x"5e",x"5b",x"5c",x"0e"),
    36 => (x"c4",x"c0",x"c0",x"c0"),
    37 => (x"4b",x"c9",x"cf",x"4c"),
    38 => (x"c9",x"e1",x"bf",x"4a"),
    39 => (x"49",x"c1",x"8a",x"71"),
    40 => (x"99",x"02",x"cf",x"87"),
    41 => (x"74",x"49",x"c1",x"84"),
    42 => (x"11",x"53",x"72",x"49"),
    43 => (x"c1",x"8a",x"71",x"99"),
    44 => (x"05",x"f1",x"87",x"c2"),
    45 => (x"87",x"26",x"4d",x"26"),
    46 => (x"4c",x"26",x"4b",x"26"),
    47 => (x"4f",x"1e",x"73",x"1e"),
    48 => (x"71",x"4b",x"e7",x"48"),
    49 => (x"c0",x"e0",x"50",x"e3"),
    50 => (x"48",x"c8",x"50",x"e3"),
    51 => (x"48",x"c6",x"50",x"e7"),
    52 => (x"48",x"c0",x"e1",x"50"),
    53 => (x"73",x"4a",x"c8",x"b7"),
    54 => (x"2a",x"c4",x"c0",x"c0"),
    55 => (x"c0",x"49",x"ca",x"81"),
    56 => (x"72",x"51",x"73",x"4a"),
    57 => (x"c3",x"ff",x"9a",x"c4"),
    58 => (x"c0",x"c0",x"c0",x"49"),
    59 => (x"cb",x"81",x"72",x"51"),
    60 => (x"e7",x"48",x"c0",x"e0"),
    61 => (x"50",x"e3",x"48",x"c8"),
    62 => (x"50",x"e3",x"48",x"c0"),
    63 => (x"50",x"e7",x"48",x"c0"),
    64 => (x"e1",x"50",x"fe",x"f4"),
    65 => (x"87",x"1e",x"73",x"1e"),
    66 => (x"c2",x"c0",x"c0",x"4b"),
    67 => (x"0f",x"fe",x"e9",x"87"),
    68 => (x"1e",x"73",x"1e",x"eb"),
    69 => (x"48",x"c3",x"ef",x"50"),
    70 => (x"e7",x"48",x"c0",x"e0"),
    71 => (x"50",x"e3",x"48",x"c8"),
    72 => (x"50",x"e3",x"48",x"c6"),
    73 => (x"50",x"e7",x"48",x"c0"),
    74 => (x"e1",x"50",x"ff",x"c2"),
    75 => (x"48",x"c1",x"9f",x"78"),
    76 => (x"e7",x"48",x"c0",x"e0"),
    77 => (x"50",x"e3",x"48",x"c4"),
    78 => (x"50",x"e3",x"48",x"c2"),
    79 => (x"50",x"e7",x"48",x"c0"),
    80 => (x"e1",x"50",x"e7",x"48"),
    81 => (x"c0",x"e0",x"50",x"e3"),
    82 => (x"48",x"c8",x"50",x"e3"),
    83 => (x"48",x"c7",x"50",x"e7"),
    84 => (x"48",x"c0",x"e1",x"50"),
    85 => (x"fc",x"f4",x"87",x"c0"),
    86 => (x"ff",x"ff",x"49",x"fd"),
    87 => (x"df",x"87",x"c0",x"fc"),
    88 => (x"c0",x"4b",x"c8",x"db"),
    89 => (x"49",x"c0",x"ed",x"f8"),
    90 => (x"87",x"cd",x"e5",x"87"),
    91 => (x"70",x"98",x"02",x"c1"),
    92 => (x"c3",x"87",x"c0",x"ff"),
    93 => (x"f0",x"4b",x"c8",x"c4"),
    94 => (x"49",x"c0",x"ed",x"e4"),
    95 => (x"87",x"d3",x"cf",x"87"),
    96 => (x"70",x"98",x"02",x"c0"),
    97 => (x"e6",x"87",x"c3",x"f0"),
    98 => (x"4b",x"c2",x"c0",x"c0"),
    99 => (x"1e",x"c7",x"c7",x"49"),
   100 => (x"c0",x"ea",x"d0",x"87"),
   101 => (x"c4",x"86",x"70",x"98"),
   102 => (x"02",x"c8",x"87",x"c3"),
   103 => (x"ff",x"4b",x"fd",x"e4"),
   104 => (x"87",x"d9",x"87",x"c7"),
   105 => (x"d3",x"49",x"c0",x"ec"),
   106 => (x"f7",x"87",x"d0",x"87"),
   107 => (x"c7",x"e8",x"49",x"c0"),
   108 => (x"ec",x"ee",x"87",x"c7"),
   109 => (x"87",x"c8",x"f1",x"49"),
   110 => (x"c0",x"ec",x"e5",x"87"),
   111 => (x"73",x"49",x"fb",x"fc"),
   112 => (x"87",x"fe",x"da",x"87"),
   113 => (x"fb",x"f2",x"87",x"38"),
   114 => (x"33",x"32",x"4f",x"53"),
   115 => (x"44",x"41",x"44",x"42"),
   116 => (x"49",x"4e",x"00",x"43"),
   117 => (x"61",x"6e",x"27",x"74"),
   118 => (x"20",x"6c",x"6f",x"61"),
   119 => (x"64",x"20",x"66",x"69"),
   120 => (x"72",x"6d",x"77",x"61"),
   121 => (x"72",x"65",x"0a",x"00"),
   122 => (x"55",x"6e",x"61",x"62"),
   123 => (x"6c",x"65",x"20",x"74"),
   124 => (x"6f",x"20",x"6c",x"6f"),
   125 => (x"63",x"61",x"74",x"65"),
   126 => (x"20",x"70",x"61",x"72"),
   127 => (x"74",x"69",x"74",x"69"),
   128 => (x"6f",x"6e",x"0a",x"00"),
   129 => (x"48",x"75",x"6e",x"74"),
   130 => (x"69",x"6e",x"67",x"20"),
   131 => (x"66",x"6f",x"72",x"20"),
   132 => (x"70",x"61",x"72",x"74"),
   133 => (x"69",x"74",x"69",x"6f"),
   134 => (x"6e",x"0a",x"00",x"49"),
   135 => (x"6e",x"69",x"74",x"69"),
   136 => (x"61",x"6c",x"69",x"7a"),
   137 => (x"69",x"6e",x"67",x"20"),
   138 => (x"53",x"44",x"20",x"63"),
   139 => (x"61",x"72",x"64",x"0a"),
   140 => (x"00",x"46",x"61",x"69"),
   141 => (x"6c",x"65",x"64",x"20"),
   142 => (x"74",x"6f",x"20",x"69"),
   143 => (x"6e",x"69",x"74",x"69"),
   144 => (x"61",x"6c",x"69",x"7a"),
   145 => (x"65",x"20",x"53",x"44"),
   146 => (x"20",x"63",x"61",x"72"),
   147 => (x"64",x"0a",x"00",x"00"),
   148 => (x"00",x"00",x"00",x"00"),
   149 => (x"00",x"00",x"08",x"33"),
   150 => (x"fc",x"0f",x"ff",x"00"),
   151 => (x"df",x"f1",x"80",x"60"),
   152 => (x"f6",x"00",x"00",x"00"),
   153 => (x"12",x"1e",x"e4",x"86"),
   154 => (x"e3",x"48",x"c3",x"ff"),
   155 => (x"50",x"e3",x"97",x"bf"),
   156 => (x"7e",x"6e",x"49",x"c3"),
   157 => (x"ff",x"99",x"e3",x"48"),
   158 => (x"c3",x"ff",x"50",x"c8"),
   159 => (x"31",x"e3",x"97",x"bf"),
   160 => (x"48",x"c8",x"a6",x"58"),
   161 => (x"c3",x"ff",x"98",x"cc"),
   162 => (x"a6",x"58",x"70",x"b1"),
   163 => (x"e3",x"48",x"c3",x"ff"),
   164 => (x"50",x"c8",x"31",x"e3"),
   165 => (x"97",x"bf",x"48",x"d0"),
   166 => (x"a6",x"58",x"c3",x"ff"),
   167 => (x"98",x"d4",x"a6",x"58"),
   168 => (x"70",x"b1",x"e3",x"48"),
   169 => (x"c3",x"ff",x"50",x"c8"),
   170 => (x"31",x"e3",x"97",x"bf"),
   171 => (x"48",x"d8",x"a6",x"58"),
   172 => (x"c3",x"ff",x"98",x"dc"),
   173 => (x"a6",x"58",x"70",x"b1"),
   174 => (x"71",x"48",x"e4",x"8e"),
   175 => (x"26",x"4f",x"0e",x"5e"),
   176 => (x"5b",x"5c",x"0e",x"1e"),
   177 => (x"71",x"4a",x"49",x"c3"),
   178 => (x"ff",x"99",x"e3",x"48"),
   179 => (x"71",x"50",x"c1",x"c0"),
   180 => (x"e4",x"bf",x"05",x"c8"),
   181 => (x"87",x"d0",x"66",x"48"),
   182 => (x"c9",x"30",x"d4",x"a6"),
   183 => (x"58",x"d0",x"66",x"49"),
   184 => (x"d8",x"29",x"c3",x"ff"),
   185 => (x"99",x"e3",x"48",x"71"),
   186 => (x"50",x"d0",x"66",x"49"),
   187 => (x"d0",x"29",x"c3",x"ff"),
   188 => (x"99",x"e3",x"48",x"71"),
   189 => (x"50",x"d0",x"66",x"49"),
   190 => (x"c8",x"29",x"c3",x"ff"),
   191 => (x"99",x"e3",x"48",x"71"),
   192 => (x"50",x"d0",x"66",x"49"),
   193 => (x"c3",x"ff",x"99",x"e3"),
   194 => (x"48",x"71",x"50",x"72"),
   195 => (x"49",x"d0",x"29",x"c3"),
   196 => (x"ff",x"99",x"e3",x"48"),
   197 => (x"71",x"50",x"e3",x"97"),
   198 => (x"bf",x"7e",x"6e",x"4b"),
   199 => (x"c3",x"ff",x"9b",x"c9"),
   200 => (x"f0",x"ff",x"4c",x"c3"),
   201 => (x"ff",x"ab",x"05",x"d9"),
   202 => (x"87",x"e3",x"48",x"c3"),
   203 => (x"ff",x"50",x"e3",x"97"),
   204 => (x"bf",x"7e",x"6e",x"4b"),
   205 => (x"c3",x"ff",x"9b",x"c1"),
   206 => (x"8c",x"02",x"c6",x"87"),
   207 => (x"c3",x"ff",x"ab",x"02"),
   208 => (x"e7",x"87",x"73",x"4a"),
   209 => (x"c4",x"b7",x"2a",x"c0"),
   210 => (x"f0",x"a2",x"49",x"c0"),
   211 => (x"e6",x"ca",x"87",x"73"),
   212 => (x"4a",x"cf",x"9a",x"c0"),
   213 => (x"f0",x"a2",x"49",x"c0"),
   214 => (x"e5",x"fe",x"87",x"73"),
   215 => (x"48",x"26",x"c2",x"87"),
   216 => (x"26",x"4d",x"26",x"4c"),
   217 => (x"26",x"4b",x"26",x"4f"),
   218 => (x"1e",x"c0",x"49",x"e3"),
   219 => (x"48",x"c3",x"ff",x"50"),
   220 => (x"c1",x"81",x"c3",x"c8"),
   221 => (x"b7",x"a9",x"04",x"f2"),
   222 => (x"87",x"26",x"4f",x"1e"),
   223 => (x"73",x"1e",x"e8",x"87"),
   224 => (x"c4",x"f8",x"df",x"4b"),
   225 => (x"c0",x"1e",x"c0",x"ff"),
   226 => (x"f0",x"c1",x"f7",x"49"),
   227 => (x"fc",x"ef",x"87",x"c4"),
   228 => (x"86",x"c1",x"a8",x"05"),
   229 => (x"c0",x"e8",x"87",x"e3"),
   230 => (x"48",x"c3",x"ff",x"50"),
   231 => (x"c1",x"c0",x"c0",x"c0"),
   232 => (x"c0",x"c0",x"1e",x"c0"),
   233 => (x"e1",x"f0",x"c1",x"e9"),
   234 => (x"49",x"fc",x"d2",x"87"),
   235 => (x"c4",x"86",x"70",x"98"),
   236 => (x"05",x"c9",x"87",x"e3"),
   237 => (x"48",x"c3",x"ff",x"50"),
   238 => (x"c1",x"48",x"cb",x"87"),
   239 => (x"fe",x"e9",x"87",x"c1"),
   240 => (x"8b",x"05",x"fe",x"ff"),
   241 => (x"87",x"c0",x"48",x"fe"),
   242 => (x"da",x"87",x"1e",x"73"),
   243 => (x"1e",x"e3",x"48",x"c3"),
   244 => (x"ff",x"50",x"d0",x"c4"),
   245 => (x"49",x"c0",x"e4",x"c8"),
   246 => (x"87",x"d3",x"4b",x"c0"),
   247 => (x"1e",x"c0",x"ff",x"f0"),
   248 => (x"c1",x"c1",x"49",x"fb"),
   249 => (x"d8",x"87",x"c4",x"86"),
   250 => (x"70",x"98",x"05",x"c9"),
   251 => (x"87",x"e3",x"48",x"c3"),
   252 => (x"ff",x"50",x"c1",x"48"),
   253 => (x"cb",x"87",x"fd",x"ef"),
   254 => (x"87",x"c1",x"8b",x"05"),
   255 => (x"ff",x"dc",x"87",x"c0"),
   256 => (x"48",x"fd",x"e0",x"87"),
   257 => (x"43",x"6d",x"64",x"5f"),
   258 => (x"69",x"6e",x"69",x"74"),
   259 => (x"0a",x"00",x"1e",x"73"),
   260 => (x"1e",x"1e",x"fd",x"d3"),
   261 => (x"87",x"c6",x"ea",x"1e"),
   262 => (x"c0",x"e1",x"f0",x"c1"),
   263 => (x"c8",x"49",x"fa",x"dd"),
   264 => (x"87",x"70",x"4b",x"1e"),
   265 => (x"d2",x"fa",x"1e",x"c0"),
   266 => (x"ed",x"fe",x"87",x"cc"),
   267 => (x"86",x"c1",x"ab",x"02"),
   268 => (x"c8",x"87",x"fe",x"d5"),
   269 => (x"87",x"c0",x"48",x"c1"),
   270 => (x"fc",x"87",x"f8",x"e8"),
   271 => (x"87",x"70",x"49",x"cf"),
   272 => (x"ff",x"ff",x"99",x"c6"),
   273 => (x"ea",x"a9",x"02",x"c8"),
   274 => (x"87",x"fd",x"fe",x"87"),
   275 => (x"c0",x"48",x"c1",x"e5"),
   276 => (x"87",x"e3",x"48",x"c3"),
   277 => (x"ff",x"50",x"c0",x"f1"),
   278 => (x"4b",x"fc",x"df",x"87"),
   279 => (x"70",x"98",x"02",x"c1"),
   280 => (x"c3",x"87",x"c0",x"1e"),
   281 => (x"c0",x"ff",x"f0",x"c1"),
   282 => (x"fa",x"49",x"f9",x"d1"),
   283 => (x"87",x"c4",x"86",x"70"),
   284 => (x"98",x"05",x"c0",x"f0"),
   285 => (x"87",x"e3",x"48",x"c3"),
   286 => (x"ff",x"50",x"e3",x"97"),
   287 => (x"bf",x"7e",x"6e",x"49"),
   288 => (x"c3",x"ff",x"99",x"e3"),
   289 => (x"48",x"c3",x"ff",x"50"),
   290 => (x"e3",x"48",x"c3",x"ff"),
   291 => (x"50",x"e3",x"48",x"c3"),
   292 => (x"ff",x"50",x"e3",x"48"),
   293 => (x"c3",x"ff",x"50",x"c1"),
   294 => (x"c0",x"99",x"02",x"c4"),
   295 => (x"87",x"c1",x"48",x"d5"),
   296 => (x"87",x"c0",x"48",x"d1"),
   297 => (x"87",x"c2",x"ab",x"05"),
   298 => (x"c4",x"87",x"c0",x"48"),
   299 => (x"c8",x"87",x"c1",x"8b"),
   300 => (x"05",x"fe",x"e5",x"87"),
   301 => (x"c0",x"48",x"26",x"fa"),
   302 => (x"ea",x"87",x"63",x"6d"),
   303 => (x"64",x"5f",x"43",x"4d"),
   304 => (x"44",x"38",x"20",x"72"),
   305 => (x"65",x"73",x"70",x"6f"),
   306 => (x"6e",x"73",x"65",x"3a"),
   307 => (x"20",x"25",x"64",x"0a"),
   308 => (x"00",x"1e",x"73",x"1e"),
   309 => (x"c1",x"c0",x"e4",x"48"),
   310 => (x"c1",x"78",x"eb",x"48"),
   311 => (x"c3",x"ef",x"50",x"c7"),
   312 => (x"4b",x"e7",x"48",x"c3"),
   313 => (x"50",x"fa",x"c0",x"87"),
   314 => (x"e7",x"48",x"c2",x"50"),
   315 => (x"e3",x"48",x"c3",x"ff"),
   316 => (x"50",x"c0",x"1e",x"c0"),
   317 => (x"e5",x"d0",x"c1",x"c0"),
   318 => (x"49",x"f7",x"c2",x"87"),
   319 => (x"c4",x"86",x"c1",x"a8"),
   320 => (x"05",x"c1",x"87",x"4b"),
   321 => (x"c2",x"ab",x"05",x"c5"),
   322 => (x"87",x"c0",x"48",x"c0"),
   323 => (x"ef",x"87",x"c1",x"8b"),
   324 => (x"05",x"ff",x"cd",x"87"),
   325 => (x"fb",x"f7",x"87",x"c1"),
   326 => (x"c0",x"e8",x"58",x"70"),
   327 => (x"98",x"05",x"cd",x"87"),
   328 => (x"c1",x"1e",x"c0",x"ff"),
   329 => (x"f0",x"c1",x"d0",x"49"),
   330 => (x"f6",x"d3",x"87",x"c4"),
   331 => (x"86",x"e3",x"48",x"c3"),
   332 => (x"ff",x"50",x"e7",x"48"),
   333 => (x"c3",x"50",x"e3",x"48"),
   334 => (x"c3",x"ff",x"50",x"c1"),
   335 => (x"48",x"f8",x"e4",x"87"),
   336 => (x"0e",x"5e",x"5b",x"5c"),
   337 => (x"5d",x"0e",x"1e",x"71"),
   338 => (x"4a",x"c0",x"4d",x"e3"),
   339 => (x"48",x"c3",x"ff",x"50"),
   340 => (x"e7",x"48",x"c2",x"50"),
   341 => (x"eb",x"48",x"c7",x"50"),
   342 => (x"e3",x"48",x"c3",x"ff"),
   343 => (x"50",x"72",x"1e",x"c0"),
   344 => (x"ff",x"f0",x"c1",x"d1"),
   345 => (x"49",x"f5",x"d6",x"87"),
   346 => (x"c4",x"86",x"70",x"98"),
   347 => (x"05",x"c1",x"c5",x"87"),
   348 => (x"c5",x"ee",x"cd",x"df"),
   349 => (x"4b",x"e3",x"48",x"c3"),
   350 => (x"ff",x"50",x"e3",x"97"),
   351 => (x"bf",x"7e",x"6e",x"49"),
   352 => (x"c3",x"ff",x"99",x"c3"),
   353 => (x"fe",x"a9",x"05",x"dd"),
   354 => (x"87",x"c0",x"4c",x"f3"),
   355 => (x"d7",x"87",x"d4",x"66"),
   356 => (x"08",x"78",x"d4",x"66"),
   357 => (x"48",x"c4",x"80",x"d8"),
   358 => (x"a6",x"58",x"c1",x"84"),
   359 => (x"c2",x"c0",x"b7",x"ac"),
   360 => (x"04",x"e8",x"87",x"c1"),
   361 => (x"4b",x"4d",x"c1",x"8b"),
   362 => (x"05",x"ff",x"c9",x"87"),
   363 => (x"e3",x"48",x"c3",x"ff"),
   364 => (x"50",x"e7",x"48",x"c3"),
   365 => (x"50",x"75",x"48",x"26"),
   366 => (x"f6",x"e5",x"87",x"1e"),
   367 => (x"73",x"1e",x"71",x"4b"),
   368 => (x"49",x"d8",x"29",x"c3"),
   369 => (x"ff",x"99",x"73",x"4a"),
   370 => (x"c8",x"2a",x"cf",x"fc"),
   371 => (x"c0",x"9a",x"72",x"b1"),
   372 => (x"73",x"4a",x"c8",x"32"),
   373 => (x"c0",x"ff",x"f0",x"c0"),
   374 => (x"c0",x"9a",x"72",x"b1"),
   375 => (x"73",x"4a",x"d8",x"32"),
   376 => (x"ff",x"c0",x"c0",x"c0"),
   377 => (x"c0",x"9a",x"72",x"b1"),
   378 => (x"71",x"48",x"c4",x"87"),
   379 => (x"26",x"4d",x"26",x"4c"),
   380 => (x"26",x"4b",x"26",x"4f"),
   381 => (x"1e",x"73",x"1e",x"71"),
   382 => (x"4b",x"49",x"c8",x"29"),
   383 => (x"c3",x"ff",x"99",x"73"),
   384 => (x"4a",x"c8",x"32",x"cf"),
   385 => (x"fc",x"c0",x"9a",x"72"),
   386 => (x"b1",x"71",x"48",x"e3"),
   387 => (x"87",x"0e",x"5e",x"5b"),
   388 => (x"5c",x"0e",x"71",x"4b"),
   389 => (x"c0",x"4c",x"d0",x"66"),
   390 => (x"48",x"c0",x"b7",x"a8"),
   391 => (x"06",x"c0",x"e3",x"87"),
   392 => (x"13",x"4a",x"cc",x"66"),
   393 => (x"97",x"bf",x"49",x"cc"),
   394 => (x"66",x"48",x"c1",x"80"),
   395 => (x"d0",x"a6",x"58",x"71"),
   396 => (x"b7",x"aa",x"02",x"c4"),
   397 => (x"87",x"c1",x"48",x"cc"),
   398 => (x"87",x"c1",x"84",x"d0"),
   399 => (x"66",x"b7",x"ac",x"04"),
   400 => (x"ff",x"dd",x"87",x"c0"),
   401 => (x"48",x"c2",x"87",x"26"),
   402 => (x"4d",x"26",x"4c",x"26"),
   403 => (x"4b",x"26",x"4f",x"0e"),
   404 => (x"5e",x"5b",x"5c",x"0e"),
   405 => (x"1e",x"c1",x"c9",x"d8"),
   406 => (x"48",x"ff",x"78",x"c1"),
   407 => (x"c8",x"f0",x"48",x"c0"),
   408 => (x"78",x"c0",x"e6",x"e9"),
   409 => (x"49",x"d9",x"f9",x"87"),
   410 => (x"c1",x"c0",x"e8",x"1e"),
   411 => (x"c0",x"49",x"fb",x"cf"),
   412 => (x"87",x"c4",x"86",x"70"),
   413 => (x"98",x"05",x"c5",x"87"),
   414 => (x"c0",x"48",x"ca",x"e5"),
   415 => (x"87",x"c0",x"4b",x"c1"),
   416 => (x"c9",x"d4",x"48",x"c1"),
   417 => (x"78",x"c8",x"1e",x"c0"),
   418 => (x"e6",x"f6",x"1e",x"c1"),
   419 => (x"c1",x"de",x"49",x"fd"),
   420 => (x"fb",x"87",x"c8",x"86"),
   421 => (x"70",x"98",x"05",x"c6"),
   422 => (x"87",x"c1",x"c9",x"d4"),
   423 => (x"48",x"c0",x"78",x"c8"),
   424 => (x"1e",x"c0",x"e6",x"ff"),
   425 => (x"1e",x"c1",x"c1",x"fa"),
   426 => (x"49",x"fd",x"e1",x"87"),
   427 => (x"c8",x"86",x"70",x"98"),
   428 => (x"05",x"c6",x"87",x"c1"),
   429 => (x"c9",x"d4",x"48",x"c0"),
   430 => (x"78",x"c8",x"1e",x"c0"),
   431 => (x"e7",x"c8",x"1e",x"c1"),
   432 => (x"c1",x"fa",x"49",x"fd"),
   433 => (x"c7",x"87",x"c8",x"86"),
   434 => (x"70",x"98",x"05",x"c5"),
   435 => (x"87",x"c0",x"48",x"c9"),
   436 => (x"d0",x"87",x"c1",x"c9"),
   437 => (x"d4",x"bf",x"1e",x"c0"),
   438 => (x"e7",x"d1",x"1e",x"c0"),
   439 => (x"e3",x"ca",x"87",x"c8"),
   440 => (x"86",x"c1",x"c9",x"d4"),
   441 => (x"bf",x"02",x"c1",x"ec"),
   442 => (x"87",x"c1",x"c0",x"e8"),
   443 => (x"4a",x"48",x"c6",x"fe"),
   444 => (x"a0",x"4c",x"c1",x"c7"),
   445 => (x"ee",x"bf",x"4b",x"c1"),
   446 => (x"c8",x"e6",x"9f",x"bf"),
   447 => (x"49",x"72",x"7e",x"c5"),
   448 => (x"d6",x"ea",x"a9",x"05"),
   449 => (x"c0",x"cc",x"87",x"c8"),
   450 => (x"a4",x"4a",x"6a",x"49"),
   451 => (x"fa",x"ec",x"87",x"70"),
   452 => (x"4b",x"db",x"87",x"c7"),
   453 => (x"fe",x"a2",x"49",x"9f"),
   454 => (x"69",x"49",x"ca",x"e9"),
   455 => (x"d5",x"a9",x"02",x"c0"),
   456 => (x"cc",x"87",x"c0",x"e4"),
   457 => (x"e6",x"49",x"d6",x"f8"),
   458 => (x"87",x"c0",x"48",x"c7"),
   459 => (x"f4",x"87",x"73",x"1e"),
   460 => (x"c0",x"e5",x"c4",x"1e"),
   461 => (x"c0",x"e1",x"f1",x"87"),
   462 => (x"c1",x"c0",x"e8",x"1e"),
   463 => (x"73",x"49",x"f7",x"ff"),
   464 => (x"87",x"cc",x"86",x"70"),
   465 => (x"98",x"05",x"c0",x"c5"),
   466 => (x"87",x"c0",x"48",x"c7"),
   467 => (x"d4",x"87",x"c0",x"e5"),
   468 => (x"dc",x"49",x"d6",x"cc"),
   469 => (x"87",x"c0",x"e7",x"e4"),
   470 => (x"1e",x"c0",x"e1",x"cc"),
   471 => (x"87",x"c8",x"1e",x"c0"),
   472 => (x"e7",x"fc",x"1e",x"c1"),
   473 => (x"c1",x"fa",x"49",x"fa"),
   474 => (x"e3",x"87",x"cc",x"86"),
   475 => (x"70",x"98",x"05",x"c0"),
   476 => (x"c9",x"87",x"c1",x"c8"),
   477 => (x"f0",x"48",x"c1",x"78"),
   478 => (x"c0",x"e4",x"87",x"c8"),
   479 => (x"1e",x"c0",x"e8",x"c5"),
   480 => (x"1e",x"c1",x"c1",x"de"),
   481 => (x"49",x"fa",x"c5",x"87"),
   482 => (x"c8",x"86",x"70",x"98"),
   483 => (x"02",x"c0",x"cf",x"87"),
   484 => (x"c0",x"e6",x"c3",x"1e"),
   485 => (x"c0",x"e0",x"d1",x"87"),
   486 => (x"c4",x"86",x"c0",x"48"),
   487 => (x"c6",x"c3",x"87",x"c1"),
   488 => (x"c8",x"e6",x"97",x"bf"),
   489 => (x"49",x"c1",x"d5",x"a9"),
   490 => (x"05",x"c0",x"cd",x"87"),
   491 => (x"c1",x"c8",x"e7",x"97"),
   492 => (x"bf",x"49",x"c2",x"ea"),
   493 => (x"a9",x"02",x"c0",x"c5"),
   494 => (x"87",x"c0",x"48",x"c5"),
   495 => (x"e4",x"87",x"c1",x"c0"),
   496 => (x"e8",x"97",x"bf",x"49"),
   497 => (x"c3",x"e9",x"a9",x"02"),
   498 => (x"c0",x"d2",x"87",x"c1"),
   499 => (x"c0",x"e8",x"97",x"bf"),
   500 => (x"49",x"c3",x"eb",x"a9"),
   501 => (x"02",x"c0",x"c5",x"87"),
   502 => (x"c0",x"48",x"c5",x"c5"),
   503 => (x"87",x"c1",x"c0",x"f3"),
   504 => (x"97",x"bf",x"49",x"99"),
   505 => (x"05",x"c0",x"cc",x"87"),
   506 => (x"c1",x"c0",x"f4",x"97"),
   507 => (x"bf",x"49",x"c2",x"a9"),
   508 => (x"02",x"c0",x"c5",x"87"),
   509 => (x"c0",x"48",x"c4",x"e9"),
   510 => (x"87",x"c1",x"c0",x"f5"),
   511 => (x"97",x"bf",x"48",x"c1"),
   512 => (x"c8",x"ec",x"58",x"c1"),
   513 => (x"88",x"c1",x"c8",x"f0"),
   514 => (x"58",x"c1",x"c0",x"f6"),
   515 => (x"97",x"bf",x"49",x"73"),
   516 => (x"81",x"c1",x"c0",x"f7"),
   517 => (x"97",x"bf",x"4a",x"c8"),
   518 => (x"32",x"c1",x"c8",x"f4"),
   519 => (x"48",x"72",x"a1",x"78"),
   520 => (x"c1",x"c0",x"f8",x"97"),
   521 => (x"bf",x"48",x"c1",x"c9"),
   522 => (x"cc",x"58",x"c1",x"c8"),
   523 => (x"f0",x"bf",x"02",x"c2"),
   524 => (x"e0",x"87",x"c8",x"1e"),
   525 => (x"c0",x"e6",x"e0",x"1e"),
   526 => (x"c1",x"c1",x"fa",x"49"),
   527 => (x"f7",x"ce",x"87",x"c8"),
   528 => (x"86",x"70",x"98",x"02"),
   529 => (x"c0",x"c5",x"87",x"c0"),
   530 => (x"48",x"c3",x"d6",x"87"),
   531 => (x"c1",x"c8",x"e8",x"bf"),
   532 => (x"48",x"c4",x"30",x"c1"),
   533 => (x"c9",x"d0",x"58",x"c1"),
   534 => (x"c8",x"e8",x"bf",x"4a"),
   535 => (x"c1",x"c9",x"c8",x"5a"),
   536 => (x"c1",x"c1",x"cd",x"97"),
   537 => (x"bf",x"49",x"c8",x"31"),
   538 => (x"c1",x"c1",x"cc",x"97"),
   539 => (x"bf",x"4b",x"a1",x"49"),
   540 => (x"c1",x"c1",x"ce",x"97"),
   541 => (x"bf",x"4b",x"d0",x"33"),
   542 => (x"73",x"a1",x"49",x"c1"),
   543 => (x"c1",x"cf",x"97",x"bf"),
   544 => (x"4b",x"d8",x"33",x"73"),
   545 => (x"a1",x"49",x"c1",x"c9"),
   546 => (x"d4",x"59",x"c1",x"c9"),
   547 => (x"c8",x"bf",x"91",x"c1"),
   548 => (x"c8",x"f4",x"bf",x"81"),
   549 => (x"c1",x"c8",x"fc",x"59"),
   550 => (x"c1",x"c1",x"d5",x"97"),
   551 => (x"bf",x"4b",x"c8",x"33"),
   552 => (x"c1",x"c1",x"d4",x"97"),
   553 => (x"bf",x"4c",x"a3",x"4b"),
   554 => (x"c1",x"c1",x"d6",x"97"),
   555 => (x"bf",x"4c",x"d0",x"34"),
   556 => (x"74",x"a3",x"4b",x"c1"),
   557 => (x"c1",x"d7",x"97",x"bf"),
   558 => (x"4c",x"cf",x"9c",x"d8"),
   559 => (x"34",x"74",x"a3",x"4b"),
   560 => (x"c1",x"c9",x"c0",x"5b"),
   561 => (x"c2",x"8b",x"73",x"92"),
   562 => (x"c1",x"c9",x"c0",x"48"),
   563 => (x"72",x"a1",x"78",x"c1"),
   564 => (x"ce",x"87",x"c1",x"c0"),
   565 => (x"fa",x"97",x"bf",x"49"),
   566 => (x"c8",x"31",x"c1",x"c0"),
   567 => (x"f9",x"97",x"bf",x"4a"),
   568 => (x"a1",x"49",x"c1",x"c9"),
   569 => (x"d0",x"59",x"c5",x"31"),
   570 => (x"c7",x"ff",x"81",x"c9"),
   571 => (x"29",x"c1",x"c9",x"c8"),
   572 => (x"59",x"c1",x"c0",x"ff"),
   573 => (x"97",x"bf",x"4a",x"c8"),
   574 => (x"32",x"c1",x"c0",x"fe"),
   575 => (x"97",x"bf",x"4b",x"a2"),
   576 => (x"4a",x"c1",x"c9",x"d4"),
   577 => (x"5a",x"c1",x"c9",x"c8"),
   578 => (x"bf",x"92",x"c1",x"c8"),
   579 => (x"f4",x"bf",x"82",x"c1"),
   580 => (x"c9",x"c4",x"5a",x"c1"),
   581 => (x"c8",x"fc",x"48",x"c0"),
   582 => (x"78",x"c1",x"c8",x"f8"),
   583 => (x"48",x"72",x"a1",x"78"),
   584 => (x"c1",x"48",x"26",x"f4"),
   585 => (x"e3",x"87",x"4e",x"6f"),
   586 => (x"20",x"70",x"61",x"72"),
   587 => (x"74",x"69",x"74",x"69"),
   588 => (x"6f",x"6e",x"20",x"73"),
   589 => (x"69",x"67",x"6e",x"61"),
   590 => (x"74",x"75",x"72",x"65"),
   591 => (x"20",x"66",x"6f",x"75"),
   592 => (x"6e",x"64",x"0a",x"00"),
   593 => (x"52",x"65",x"61",x"64"),
   594 => (x"69",x"6e",x"67",x"20"),
   595 => (x"62",x"6f",x"6f",x"74"),
   596 => (x"20",x"73",x"65",x"63"),
   597 => (x"74",x"6f",x"72",x"20"),
   598 => (x"25",x"64",x"0a",x"00"),
   599 => (x"52",x"65",x"61",x"64"),
   600 => (x"20",x"62",x"6f",x"6f"),
   601 => (x"74",x"20",x"73",x"65"),
   602 => (x"63",x"74",x"6f",x"72"),
   603 => (x"20",x"66",x"72",x"6f"),
   604 => (x"6d",x"20",x"66",x"69"),
   605 => (x"72",x"73",x"74",x"20"),
   606 => (x"70",x"61",x"72",x"74"),
   607 => (x"69",x"74",x"69",x"6f"),
   608 => (x"6e",x"0a",x"00",x"55"),
   609 => (x"6e",x"73",x"75",x"70"),
   610 => (x"70",x"6f",x"72",x"74"),
   611 => (x"65",x"64",x"20",x"70"),
   612 => (x"61",x"72",x"74",x"69"),
   613 => (x"74",x"69",x"6f",x"6e"),
   614 => (x"20",x"74",x"79",x"70"),
   615 => (x"65",x"21",x"0d",x"00"),
   616 => (x"46",x"41",x"54",x"33"),
   617 => (x"32",x"20",x"20",x"20"),
   618 => (x"00",x"52",x"65",x"61"),
   619 => (x"64",x"69",x"6e",x"67"),
   620 => (x"20",x"4d",x"42",x"52"),
   621 => (x"0a",x"00",x"46",x"41"),
   622 => (x"54",x"31",x"36",x"20"),
   623 => (x"20",x"20",x"00",x"46"),
   624 => (x"41",x"54",x"33",x"32"),
   625 => (x"20",x"20",x"20",x"00"),
   626 => (x"46",x"41",x"54",x"31"),
   627 => (x"32",x"20",x"20",x"20"),
   628 => (x"00",x"50",x"61",x"72"),
   629 => (x"74",x"69",x"74",x"69"),
   630 => (x"6f",x"6e",x"63",x"6f"),
   631 => (x"75",x"6e",x"74",x"20"),
   632 => (x"25",x"64",x"0a",x"00"),
   633 => (x"48",x"75",x"6e",x"74"),
   634 => (x"69",x"6e",x"67",x"20"),
   635 => (x"66",x"6f",x"72",x"20"),
   636 => (x"66",x"69",x"6c",x"65"),
   637 => (x"73",x"79",x"73",x"74"),
   638 => (x"65",x"6d",x"0a",x"00"),
   639 => (x"46",x"41",x"54",x"33"),
   640 => (x"32",x"20",x"20",x"20"),
   641 => (x"00",x"46",x"41",x"54"),
   642 => (x"31",x"36",x"20",x"20"),
   643 => (x"20",x"00",x"0e",x"5e"),
   644 => (x"5b",x"5c",x"5d",x"0e"),
   645 => (x"71",x"4a",x"c1",x"c8"),
   646 => (x"f0",x"bf",x"02",x"cc"),
   647 => (x"87",x"72",x"4b",x"c7"),
   648 => (x"b7",x"2b",x"72",x"4c"),
   649 => (x"c1",x"ff",x"9c",x"ca"),
   650 => (x"87",x"72",x"4b",x"c8"),
   651 => (x"b7",x"2b",x"72",x"4c"),
   652 => (x"c3",x"ff",x"9c",x"c1"),
   653 => (x"c9",x"d8",x"bf",x"ab"),
   654 => (x"02",x"de",x"87",x"c1"),
   655 => (x"c0",x"e8",x"1e",x"c1"),
   656 => (x"c8",x"f4",x"bf",x"49"),
   657 => (x"73",x"81",x"eb",x"f7"),
   658 => (x"87",x"c4",x"86",x"70"),
   659 => (x"98",x"05",x"c5",x"87"),
   660 => (x"c0",x"48",x"c0",x"f5"),
   661 => (x"87",x"c1",x"c9",x"dc"),
   662 => (x"5b",x"c1",x"c8",x"f0"),
   663 => (x"bf",x"02",x"d8",x"87"),
   664 => (x"74",x"4a",x"c4",x"92"),
   665 => (x"c1",x"c0",x"e8",x"82"),
   666 => (x"6a",x"49",x"ed",x"ce"),
   667 => (x"87",x"70",x"49",x"4d"),
   668 => (x"cf",x"ff",x"ff",x"ff"),
   669 => (x"ff",x"9d",x"d0",x"87"),
   670 => (x"74",x"4a",x"c2",x"92"),
   671 => (x"c1",x"c0",x"e8",x"82"),
   672 => (x"9f",x"6a",x"49",x"ed"),
   673 => (x"ee",x"87",x"70",x"4d"),
   674 => (x"75",x"48",x"ee",x"fa"),
   675 => (x"87",x"0e",x"5e",x"5b"),
   676 => (x"5c",x"5d",x"0e",x"f4"),
   677 => (x"86",x"71",x"4c",x"c0"),
   678 => (x"4b",x"c1",x"c9",x"d8"),
   679 => (x"48",x"ff",x"78",x"c1"),
   680 => (x"c8",x"fc",x"bf",x"4d"),
   681 => (x"c1",x"c9",x"c0",x"bf"),
   682 => (x"7e",x"c1",x"c8",x"f0"),
   683 => (x"bf",x"02",x"c9",x"87"),
   684 => (x"c1",x"c8",x"e8",x"bf"),
   685 => (x"4a",x"c4",x"32",x"c7"),
   686 => (x"87",x"c1",x"c9",x"c4"),
   687 => (x"bf",x"4a",x"c4",x"32"),
   688 => (x"c8",x"a6",x"5a",x"c8"),
   689 => (x"a6",x"48",x"c0",x"78"),
   690 => (x"c4",x"66",x"48",x"c0"),
   691 => (x"a8",x"06",x"c3",x"cc"),
   692 => (x"87",x"c8",x"66",x"49"),
   693 => (x"cf",x"99",x"05",x"c0"),
   694 => (x"e2",x"87",x"6e",x"1e"),
   695 => (x"c0",x"ef",x"de",x"1e"),
   696 => (x"d3",x"c6",x"87",x"c1"),
   697 => (x"c0",x"e8",x"1e",x"cc"),
   698 => (x"66",x"49",x"48",x"c1"),
   699 => (x"80",x"d0",x"a6",x"58"),
   700 => (x"71",x"e9",x"cc",x"87"),
   701 => (x"cc",x"86",x"c1",x"c0"),
   702 => (x"e8",x"4b",x"c3",x"87"),
   703 => (x"c0",x"e0",x"83",x"97"),
   704 => (x"6b",x"49",x"99",x"02"),
   705 => (x"c2",x"c4",x"87",x"97"),
   706 => (x"6b",x"49",x"c3",x"e5"),
   707 => (x"a9",x"02",x"c1",x"fa"),
   708 => (x"87",x"cb",x"a3",x"49"),
   709 => (x"97",x"69",x"49",x"d8"),
   710 => (x"99",x"05",x"c1",x"ee"),
   711 => (x"87",x"cb",x"1e",x"c0"),
   712 => (x"e0",x"66",x"1e",x"73"),
   713 => (x"49",x"eb",x"e5",x"87"),
   714 => (x"c8",x"86",x"70",x"98"),
   715 => (x"05",x"c1",x"db",x"87"),
   716 => (x"dc",x"a3",x"4a",x"6a"),
   717 => (x"49",x"ea",x"c3",x"87"),
   718 => (x"70",x"4a",x"c4",x"a4"),
   719 => (x"49",x"72",x"79",x"da"),
   720 => (x"a3",x"4a",x"9f",x"6a"),
   721 => (x"49",x"ea",x"ec",x"87"),
   722 => (x"70",x"7e",x"c1",x"c8"),
   723 => (x"f0",x"bf",x"02",x"d8"),
   724 => (x"87",x"d4",x"a3",x"4a"),
   725 => (x"9f",x"6a",x"49",x"ea"),
   726 => (x"da",x"87",x"70",x"49"),
   727 => (x"c0",x"ff",x"ff",x"99"),
   728 => (x"71",x"48",x"d0",x"30"),
   729 => (x"c8",x"a6",x"58",x"c5"),
   730 => (x"87",x"c4",x"a6",x"48"),
   731 => (x"c0",x"78",x"c4",x"66"),
   732 => (x"4a",x"6e",x"82",x"c8"),
   733 => (x"a4",x"49",x"72",x"79"),
   734 => (x"c0",x"7c",x"dc",x"66"),
   735 => (x"1e",x"c0",x"ef",x"fb"),
   736 => (x"1e",x"d0",x"e5",x"87"),
   737 => (x"c8",x"86",x"c1",x"48"),
   738 => (x"c1",x"ce",x"87",x"c8"),
   739 => (x"66",x"48",x"c1",x"80"),
   740 => (x"cc",x"a6",x"58",x"c8"),
   741 => (x"66",x"48",x"c4",x"66"),
   742 => (x"a8",x"04",x"fc",x"f4"),
   743 => (x"87",x"c1",x"c8",x"f0"),
   744 => (x"bf",x"02",x"c0",x"f2"),
   745 => (x"87",x"75",x"49",x"f9"),
   746 => (x"e4",x"87",x"70",x"4d"),
   747 => (x"1e",x"c0",x"f0",x"cc"),
   748 => (x"1e",x"cf",x"f5",x"87"),
   749 => (x"c8",x"86",x"75",x"49"),
   750 => (x"cf",x"ff",x"ff",x"ff"),
   751 => (x"f8",x"99",x"a9",x"02"),
   752 => (x"d5",x"87",x"75",x"49"),
   753 => (x"c2",x"89",x"c1",x"c8"),
   754 => (x"e8",x"bf",x"91",x"c1"),
   755 => (x"c8",x"f8",x"bf",x"48"),
   756 => (x"71",x"80",x"70",x"7e"),
   757 => (x"fb",x"ec",x"87",x"c0"),
   758 => (x"48",x"f4",x"8e",x"e9"),
   759 => (x"e9",x"87",x"52",x"65"),
   760 => (x"61",x"64",x"69",x"6e"),
   761 => (x"67",x"20",x"64",x"69"),
   762 => (x"72",x"65",x"63",x"74"),
   763 => (x"6f",x"72",x"79",x"20"),
   764 => (x"73",x"65",x"63",x"74"),
   765 => (x"6f",x"72",x"20",x"25"),
   766 => (x"64",x"0a",x"00",x"66"),
   767 => (x"69",x"6c",x"65",x"20"),
   768 => (x"22",x"25",x"73",x"22"),
   769 => (x"20",x"66",x"6f",x"75"),
   770 => (x"6e",x"64",x"0d",x"00"),
   771 => (x"47",x"65",x"74",x"46"),
   772 => (x"41",x"54",x"4c",x"69"),
   773 => (x"6e",x"6b",x"20",x"72"),
   774 => (x"65",x"74",x"75",x"72"),
   775 => (x"6e",x"65",x"64",x"20"),
   776 => (x"25",x"64",x"0a",x"00"),
   777 => (x"0e",x"5e",x"5b",x"5c"),
   778 => (x"5d",x"0e",x"1e",x"71"),
   779 => (x"4b",x"1e",x"c1",x"c9"),
   780 => (x"dc",x"49",x"f9",x"d8"),
   781 => (x"87",x"c4",x"86",x"70"),
   782 => (x"98",x"02",x"c1",x"f5"),
   783 => (x"87",x"c1",x"c9",x"e0"),
   784 => (x"bf",x"49",x"c7",x"ff"),
   785 => (x"81",x"c9",x"29",x"71"),
   786 => (x"7e",x"c0",x"4d",x"4c"),
   787 => (x"6e",x"48",x"c0",x"b7"),
   788 => (x"a8",x"06",x"c1",x"ec"),
   789 => (x"87",x"c1",x"c8",x"f8"),
   790 => (x"bf",x"49",x"c1",x"c9"),
   791 => (x"e4",x"bf",x"4a",x"c2"),
   792 => (x"8a",x"c1",x"c8",x"e8"),
   793 => (x"bf",x"92",x"72",x"a1"),
   794 => (x"49",x"c1",x"c8",x"ec"),
   795 => (x"bf",x"4a",x"74",x"9a"),
   796 => (x"72",x"a1",x"49",x"d4"),
   797 => (x"66",x"1e",x"71",x"e3"),
   798 => (x"c6",x"87",x"c4",x"86"),
   799 => (x"70",x"98",x"05",x"c5"),
   800 => (x"87",x"c0",x"48",x"c1"),
   801 => (x"c0",x"87",x"c1",x"84"),
   802 => (x"c1",x"c8",x"ec",x"bf"),
   803 => (x"49",x"74",x"99",x"05"),
   804 => (x"cc",x"87",x"c1",x"c9"),
   805 => (x"e4",x"bf",x"49",x"f5"),
   806 => (x"f4",x"87",x"c1",x"c9"),
   807 => (x"e8",x"58",x"d4",x"66"),
   808 => (x"48",x"c8",x"c0",x"80"),
   809 => (x"d8",x"a6",x"58",x"c1"),
   810 => (x"85",x"6e",x"b7",x"ad"),
   811 => (x"04",x"fe",x"e5",x"87"),
   812 => (x"cf",x"87",x"73",x"1e"),
   813 => (x"c0",x"f3",x"ca",x"1e"),
   814 => (x"cb",x"ee",x"87",x"c8"),
   815 => (x"86",x"c0",x"48",x"c5"),
   816 => (x"87",x"c1",x"c9",x"e0"),
   817 => (x"bf",x"48",x"26",x"e5"),
   818 => (x"fd",x"87",x"43",x"61"),
   819 => (x"6e",x"27",x"74",x"20"),
   820 => (x"6f",x"70",x"65",x"6e"),
   821 => (x"20",x"25",x"73",x"0a"),
   822 => (x"00",x"1e",x"f3",x"48"),
   823 => (x"71",x"50",x"48",x"26"),
   824 => (x"4f",x"0e",x"5e",x"5b"),
   825 => (x"5c",x"0e",x"71",x"4b"),
   826 => (x"c0",x"4c",x"13",x"4a"),
   827 => (x"9a",x"02",x"cc",x"87"),
   828 => (x"72",x"49",x"e5",x"87"),
   829 => (x"c1",x"84",x"13",x"4a"),
   830 => (x"9a",x"05",x"f4",x"87"),
   831 => (x"74",x"48",x"c2",x"87"),
   832 => (x"26",x"4d",x"26",x"4c"),
   833 => (x"26",x"4b",x"26",x"4f"),
   834 => (x"0e",x"5e",x"5b",x"5c"),
   835 => (x"5d",x"0e",x"fc",x"86"),
   836 => (x"71",x"4a",x"c0",x"e0"),
   837 => (x"66",x"4c",x"d5",x"cf"),
   838 => (x"a7",x"4b",x"c0",x"7e"),
   839 => (x"72",x"9a",x"05",x"ce"),
   840 => (x"87",x"d5",x"c5",x"a7"),
   841 => (x"4b",x"d5",x"c0",x"a7"),
   842 => (x"48",x"c0",x"f0",x"50"),
   843 => (x"c1",x"c9",x"87",x"72"),
   844 => (x"9a",x"02",x"c0",x"e5"),
   845 => (x"87",x"d4",x"66",x"4d"),
   846 => (x"72",x"1e",x"72",x"49"),
   847 => (x"75",x"4a",x"c9",x"fc"),
   848 => (x"87",x"26",x"4a",x"c1"),
   849 => (x"e2",x"a7",x"81",x"11"),
   850 => (x"53",x"72",x"49",x"75"),
   851 => (x"4a",x"c9",x"ed",x"87"),
   852 => (x"70",x"4a",x"c1",x"8c"),
   853 => (x"72",x"9a",x"05",x"ff"),
   854 => (x"de",x"87",x"c0",x"b7"),
   855 => (x"ac",x"06",x"d8",x"87"),
   856 => (x"c0",x"e4",x"66",x"02"),
   857 => (x"c5",x"87",x"c0",x"f0"),
   858 => (x"4a",x"c3",x"87",x"c0"),
   859 => (x"e0",x"4a",x"72",x"53"),
   860 => (x"c1",x"8c",x"c0",x"b7"),
   861 => (x"ac",x"01",x"e8",x"87"),
   862 => (x"d3",x"ed",x"a7",x"ab"),
   863 => (x"02",x"dd",x"87",x"d8"),
   864 => (x"66",x"4c",x"dc",x"66"),
   865 => (x"1e",x"c1",x"8b",x"97"),
   866 => (x"6b",x"49",x"74",x"0f"),
   867 => (x"c4",x"86",x"6e",x"48"),
   868 => (x"c1",x"80",x"70",x"7e"),
   869 => (x"d3",x"d1",x"a7",x"ab"),
   870 => (x"05",x"ff",x"e6",x"87"),
   871 => (x"6e",x"48",x"fc",x"8e"),
   872 => (x"26",x"4d",x"26",x"4c"),
   873 => (x"26",x"4b",x"26",x"4f"),
   874 => (x"30",x"31",x"32",x"33"),
   875 => (x"34",x"35",x"36",x"37"),
   876 => (x"38",x"39",x"41",x"42"),
   877 => (x"43",x"44",x"45",x"46"),
   878 => (x"00",x"0e",x"5e",x"5b"),
   879 => (x"5c",x"5d",x"0e",x"71"),
   880 => (x"4b",x"ff",x"4d",x"13"),
   881 => (x"4c",x"9c",x"02",x"d7"),
   882 => (x"87",x"c1",x"85",x"d4"),
   883 => (x"66",x"1e",x"74",x"49"),
   884 => (x"d4",x"66",x"0f",x"c4"),
   885 => (x"86",x"74",x"a8",x"05"),
   886 => (x"c6",x"87",x"13",x"4c"),
   887 => (x"9c",x"05",x"e9",x"87"),
   888 => (x"75",x"48",x"26",x"4d"),
   889 => (x"26",x"4c",x"26",x"4b"),
   890 => (x"26",x"4f",x"0e",x"5e"),
   891 => (x"5b",x"5c",x"5d",x"0e"),
   892 => (x"e8",x"86",x"71",x"7e"),
   893 => (x"c0",x"e8",x"66",x"4d"),
   894 => (x"c0",x"4c",x"c8",x"a6"),
   895 => (x"48",x"c0",x"78",x"6e"),
   896 => (x"97",x"bf",x"4b",x"6e"),
   897 => (x"48",x"c1",x"80",x"70"),
   898 => (x"7e",x"73",x"9b",x"02"),
   899 => (x"c6",x"ce",x"87",x"c8"),
   900 => (x"66",x"02",x"c5",x"d7"),
   901 => (x"87",x"cc",x"a6",x"48"),
   902 => (x"c0",x"78",x"fc",x"80"),
   903 => (x"c0",x"78",x"73",x"4a"),
   904 => (x"c0",x"e0",x"8a",x"02"),
   905 => (x"c3",x"c2",x"87",x"c3"),
   906 => (x"8a",x"02",x"c2",x"fc"),
   907 => (x"87",x"c2",x"8a",x"02"),
   908 => (x"c2",x"e4",x"87",x"8a"),
   909 => (x"02",x"c2",x"f1",x"87"),
   910 => (x"c4",x"8a",x"02",x"c2"),
   911 => (x"eb",x"87",x"c2",x"8a"),
   912 => (x"02",x"c2",x"e5",x"87"),
   913 => (x"c3",x"8a",x"02",x"c2"),
   914 => (x"e7",x"87",x"d4",x"8a"),
   915 => (x"02",x"c0",x"f4",x"87"),
   916 => (x"8a",x"02",x"c0",x"ff"),
   917 => (x"87",x"ca",x"8a",x"02"),
   918 => (x"c0",x"f1",x"87",x"c1"),
   919 => (x"8a",x"02",x"c1",x"df"),
   920 => (x"87",x"8a",x"02",x"df"),
   921 => (x"87",x"c8",x"8a",x"02"),
   922 => (x"c1",x"cd",x"87",x"c4"),
   923 => (x"8a",x"02",x"c0",x"e3"),
   924 => (x"87",x"c3",x"8a",x"02"),
   925 => (x"c0",x"e5",x"87",x"c2"),
   926 => (x"8a",x"02",x"c8",x"87"),
   927 => (x"c3",x"8a",x"02",x"d3"),
   928 => (x"87",x"c1",x"f9",x"87"),
   929 => (x"cc",x"a6",x"48",x"ca"),
   930 => (x"78",x"c2",x"d2",x"87"),
   931 => (x"cc",x"a6",x"48",x"c2"),
   932 => (x"78",x"c2",x"ca",x"87"),
   933 => (x"cc",x"a6",x"48",x"d0"),
   934 => (x"78",x"c2",x"c2",x"87"),
   935 => (x"c0",x"f0",x"66",x"1e"),
   936 => (x"c0",x"f0",x"66",x"1e"),
   937 => (x"c4",x"85",x"75",x"4a"),
   938 => (x"c4",x"8a",x"6a",x"49"),
   939 => (x"fc",x"ca",x"87",x"c8"),
   940 => (x"86",x"70",x"49",x"a4"),
   941 => (x"4c",x"c1",x"e6",x"87"),
   942 => (x"c8",x"a6",x"48",x"c1"),
   943 => (x"78",x"c1",x"de",x"87"),
   944 => (x"c0",x"f0",x"66",x"1e"),
   945 => (x"c4",x"85",x"75",x"4a"),
   946 => (x"c4",x"8a",x"6a",x"49"),
   947 => (x"c0",x"f0",x"66",x"0f"),
   948 => (x"c4",x"86",x"c1",x"84"),
   949 => (x"c1",x"c7",x"87",x"c0"),
   950 => (x"f0",x"66",x"1e",x"c0"),
   951 => (x"e5",x"49",x"c0",x"f0"),
   952 => (x"66",x"0f",x"c4",x"86"),
   953 => (x"c1",x"84",x"c0",x"f5"),
   954 => (x"87",x"c8",x"a6",x"48"),
   955 => (x"c1",x"78",x"c0",x"ed"),
   956 => (x"87",x"d0",x"a6",x"48"),
   957 => (x"c1",x"78",x"f8",x"80"),
   958 => (x"c1",x"78",x"c0",x"e1"),
   959 => (x"87",x"c0",x"f0",x"ab"),
   960 => (x"06",x"db",x"87",x"c0"),
   961 => (x"f9",x"ab",x"03",x"d5"),
   962 => (x"87",x"d4",x"66",x"49"),
   963 => (x"ca",x"91",x"73",x"4a"),
   964 => (x"c0",x"f0",x"8a",x"d4"),
   965 => (x"a6",x"48",x"72",x"a1"),
   966 => (x"78",x"c8",x"a6",x"48"),
   967 => (x"c1",x"78",x"cc",x"66"),
   968 => (x"02",x"c1",x"e9",x"87"),
   969 => (x"c4",x"85",x"75",x"49"),
   970 => (x"c4",x"89",x"a6",x"48"),
   971 => (x"69",x"78",x"c1",x"e4"),
   972 => (x"ab",x"05",x"d8",x"87"),
   973 => (x"c4",x"66",x"48",x"c0"),
   974 => (x"b7",x"a8",x"03",x"cf"),
   975 => (x"87",x"c0",x"ed",x"49"),
   976 => (x"f6",x"d6",x"87",x"c4"),
   977 => (x"66",x"48",x"c0",x"08"),
   978 => (x"88",x"c8",x"a6",x"58"),
   979 => (x"d0",x"66",x"1e",x"d8"),
   980 => (x"66",x"1e",x"c0",x"f8"),
   981 => (x"66",x"1e",x"c0",x"f8"),
   982 => (x"66",x"1e",x"dc",x"66"),
   983 => (x"1e",x"d8",x"66",x"49"),
   984 => (x"f6",x"e5",x"87",x"d4"),
   985 => (x"86",x"70",x"49",x"a4"),
   986 => (x"4c",x"c0",x"e1",x"87"),
   987 => (x"c0",x"e5",x"ab",x"05"),
   988 => (x"cf",x"87",x"d0",x"a6"),
   989 => (x"48",x"c0",x"78",x"c4"),
   990 => (x"80",x"c0",x"78",x"f4"),
   991 => (x"80",x"c1",x"78",x"cc"),
   992 => (x"87",x"c0",x"f0",x"66"),
   993 => (x"1e",x"73",x"49",x"c0"),
   994 => (x"f0",x"66",x"0f",x"c4"),
   995 => (x"86",x"6e",x"97",x"bf"),
   996 => (x"4b",x"6e",x"48",x"c1"),
   997 => (x"80",x"70",x"7e",x"73"),
   998 => (x"9b",x"05",x"f9",x"f2"),
   999 => (x"87",x"74",x"48",x"e8"),
  1000 => (x"8e",x"26",x"4d",x"26"),
  1001 => (x"4c",x"26",x"4b",x"26"),
  1002 => (x"4f",x"1e",x"c0",x"1e"),
  1003 => (x"f4",x"ea",x"a7",x"1e"),
  1004 => (x"d0",x"a6",x"1e",x"d0"),
  1005 => (x"66",x"49",x"f8",x"f1"),
  1006 => (x"87",x"f4",x"8e",x"26"),
  1007 => (x"4f",x"1e",x"73",x"1e"),
  1008 => (x"72",x"9a",x"02",x"c0"),
  1009 => (x"e7",x"87",x"c0",x"48"),
  1010 => (x"c1",x"4b",x"72",x"a9"),
  1011 => (x"06",x"d1",x"87",x"72"),
  1012 => (x"82",x"06",x"c9",x"87"),
  1013 => (x"73",x"83",x"72",x"a9"),
  1014 => (x"01",x"f4",x"87",x"c3"),
  1015 => (x"87",x"c1",x"b2",x"3a"),
  1016 => (x"72",x"a9",x"03",x"89"),
  1017 => (x"73",x"80",x"07",x"c1"),
  1018 => (x"2a",x"2b",x"05",x"f3"),
  1019 => (x"87",x"26",x"4b",x"26"),
  1020 => (x"4f",x"1e",x"75",x"1e"),
  1021 => (x"c4",x"4d",x"71",x"b7"),
  1022 => (x"a1",x"04",x"ff",x"b9"),
  1023 => (x"c1",x"81",x"c3",x"bd"),
  1024 => (x"07",x"72",x"b7",x"a2"),
  1025 => (x"04",x"ff",x"ba",x"c1"),
  1026 => (x"82",x"c1",x"bd",x"07"),
  1027 => (x"fe",x"ee",x"87",x"c1"),
  1028 => (x"2d",x"04",x"ff",x"b8"),
  1029 => (x"c1",x"80",x"07",x"2d"),
  1030 => (x"04",x"ff",x"b9",x"c1"),
  1031 => (x"81",x"07",x"26",x"4d"),
  1032 => (x"26",x"4f",x"26",x"4d"),
	others => (others => x"00")
);

-- Xilinx XST attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "no_rw_check";

-- Altera Quartus attributes
attribute ramstyle: string;
attribute ramstyle of ram: signal is "no_rw_check";

signal q_local : word_t;
signal q2_local : word_t;

begin
    
	process(clk,q_local)
	begin

		q(31 downto 24)<=q_local(0);
		q(23 downto 16)<=q_local(1);
		q(15 downto 8)<=q_local(2);
		q(7 downto 0)<=q_local(3);

		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel(3) = '1') then
					ram(to_integer(unsigned(addr)))(3) <= d(7 downto 0);
				end if;
				if bytesel(2) = '1' then
					ram(to_integer(unsigned(addr)))(2) <= d(15 downto 8);
				end if;
				if bytesel(1) = '1' then
					ram(to_integer(unsigned(addr)))(1) <= d(23 downto 16);
				end if;
				if bytesel(0) = '1' then
					ram(to_integer(unsigned(addr)))(0) <= d(31 downto 24);
				end if;
			end if;
			q_local <= ram(to_integer(unsigned(addr)));
		end if;
	end process;

	-- Second port
	
	process(clk,q2_local)
	begin

		q2(31 downto 24)<=q2_local(0);
		q2(23 downto 16)<=q2_local(1);
		q2(15 downto 8)<=q2_local(2);
		q2(7 downto 0)<=q2_local(3);

		if(rising_edge(clk)) then 
			if(we2 = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel2(3) = '1') then
					ram(to_integer(unsigned(addr2)))(3) <= d2(7 downto 0);
				end if;
				if bytesel2(2) = '1' then
					ram(to_integer(unsigned(addr2)))(2) <= d2(15 downto 8);
				end if;
				if bytesel2(1) = '1' then
					ram(to_integer(unsigned(addr2)))(1) <= d2(23 downto 16);
				end if;
				if bytesel2(0) = '1' then
					ram(to_integer(unsigned(addr2)))(0) <= d2(31 downto 24);
				end if;
			end if;
			q2_local <= ram(to_integer(unsigned(addr2)));
		end if;
	end process;

end arch;

