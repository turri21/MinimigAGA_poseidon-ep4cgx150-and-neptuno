library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM-2 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
type ram_type is array (0 to 2 ** (maxAddrBitBRAM-3) - 1) of word_t;

signal ram : ram_type :=
(
     0 => (x"01",x"da",x"87",x"04"),
     1 => (x"dd",x"87",x"0e",x"58"),
     2 => (x"5e",x"59",x"5a",x"0e"),
     3 => (x"27",x"00",x"00",x"00"),
     4 => (x"2c",x"0f",x"26",x"4a"),
     5 => (x"26",x"49",x"26",x"48"),
     6 => (x"ff",x"80",x"26",x"08"),
     7 => (x"4f",x"27",x"00",x"00"),
     8 => (x"00",x"2d",x"4f",x"27"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"4f",x"00",x"fd",x"87"),
    11 => (x"4f",x"c1",x"ce",x"c4"),
    12 => (x"4e",x"c9",x"c0",x"86"),
    13 => (x"c1",x"ce",x"c4",x"49"),
    14 => (x"c1",x"c4",x"e0",x"48"),
    15 => (x"89",x"d0",x"89",x"03"),
    16 => (x"c0",x"40",x"40",x"40"),
    17 => (x"40",x"f6",x"87",x"d0"),
    18 => (x"81",x"05",x"c0",x"50"),
    19 => (x"c1",x"89",x"05",x"f9"),
    20 => (x"87",x"c1",x"c4",x"e0"),
    21 => (x"4d",x"c1",x"c4",x"e0"),
    22 => (x"4c",x"74",x"ad",x"02"),
    23 => (x"c4",x"87",x"24",x"0f"),
    24 => (x"f7",x"87",x"c2",x"e1"),
    25 => (x"87",x"c1",x"c4",x"e0"),
    26 => (x"4d",x"c1",x"c4",x"e0"),
    27 => (x"4c",x"74",x"ad",x"02"),
    28 => (x"c6",x"87",x"c4",x"8c"),
    29 => (x"6c",x"0f",x"f5",x"87"),
    30 => (x"00",x"fd",x"87",x"0e"),
    31 => (x"5e",x"5b",x"5c",x"0e"),
    32 => (x"c8",x"c0",x"c0",x"c0"),
    33 => (x"4b",x"c9",x"c5",x"4c"),
    34 => (x"c9",x"d7",x"bf",x"4a"),
    35 => (x"72",x"49",x"c1",x"8a"),
    36 => (x"71",x"99",x"02",x"cf"),
    37 => (x"87",x"74",x"49",x"c1"),
    38 => (x"84",x"11",x"53",x"72"),
    39 => (x"49",x"c1",x"8a",x"71"),
    40 => (x"99",x"05",x"f1",x"87"),
    41 => (x"c2",x"87",x"26",x"4d"),
    42 => (x"26",x"4c",x"26",x"4b"),
    43 => (x"26",x"4f",x"1e",x"73"),
    44 => (x"1e",x"71",x"4b",x"e7"),
    45 => (x"48",x"c0",x"e0",x"50"),
    46 => (x"e3",x"48",x"c8",x"50"),
    47 => (x"e3",x"48",x"c6",x"50"),
    48 => (x"e7",x"48",x"c0",x"e1"),
    49 => (x"50",x"73",x"4a",x"c8"),
    50 => (x"b7",x"2a",x"c8",x"c0"),
    51 => (x"c0",x"c0",x"49",x"ca"),
    52 => (x"81",x"71",x"0a",x"97"),
    53 => (x"7a",x"73",x"4a",x"c3"),
    54 => (x"ff",x"9a",x"c8",x"c0"),
    55 => (x"c0",x"c0",x"49",x"cb"),
    56 => (x"81",x"71",x"0a",x"97"),
    57 => (x"7a",x"e7",x"48",x"c0"),
    58 => (x"e0",x"50",x"e3",x"48"),
    59 => (x"c8",x"50",x"e3",x"48"),
    60 => (x"c0",x"50",x"e7",x"48"),
    61 => (x"c0",x"e1",x"50",x"fe"),
    62 => (x"f0",x"87",x"1e",x"73"),
    63 => (x"1e",x"c2",x"c0",x"c0"),
    64 => (x"4b",x"73",x"0f",x"fe"),
    65 => (x"e4",x"87",x"1e",x"73"),
    66 => (x"1e",x"eb",x"48",x"c3"),
    67 => (x"ef",x"50",x"e7",x"48"),
    68 => (x"c0",x"e0",x"50",x"e3"),
    69 => (x"48",x"c8",x"50",x"e3"),
    70 => (x"48",x"c6",x"50",x"e7"),
    71 => (x"48",x"c0",x"e1",x"50"),
    72 => (x"ff",x"c2",x"48",x"c1"),
    73 => (x"9f",x"78",x"e7",x"48"),
    74 => (x"c0",x"e0",x"50",x"e3"),
    75 => (x"48",x"c4",x"50",x"e3"),
    76 => (x"48",x"c2",x"50",x"e7"),
    77 => (x"48",x"c0",x"e1",x"50"),
    78 => (x"e7",x"48",x"c0",x"e0"),
    79 => (x"50",x"e3",x"48",x"c8"),
    80 => (x"50",x"e3",x"48",x"c7"),
    81 => (x"50",x"e7",x"48",x"c0"),
    82 => (x"e1",x"50",x"fc",x"ee"),
    83 => (x"87",x"c0",x"ff",x"ff"),
    84 => (x"49",x"fd",x"da",x"87"),
    85 => (x"c0",x"fc",x"c0",x"4b"),
    86 => (x"c8",x"d1",x"49",x"c0"),
    87 => (x"f1",x"eb",x"87",x"d0"),
    88 => (x"f9",x"87",x"70",x"98"),
    89 => (x"02",x"c1",x"c3",x"87"),
    90 => (x"c0",x"ff",x"f0",x"4b"),
    91 => (x"c7",x"fa",x"49",x"c0"),
    92 => (x"f1",x"d7",x"87",x"d6"),
    93 => (x"ec",x"87",x"70",x"98"),
    94 => (x"02",x"c0",x"e6",x"87"),
    95 => (x"c3",x"f0",x"4b",x"c2"),
    96 => (x"c0",x"c0",x"1e",x"c6"),
    97 => (x"fd",x"49",x"c0",x"ee"),
    98 => (x"cd",x"87",x"c4",x"86"),
    99 => (x"70",x"98",x"02",x"c8"),
   100 => (x"87",x"c3",x"ff",x"4b"),
   101 => (x"fd",x"e3",x"87",x"d9"),
   102 => (x"87",x"c7",x"c9",x"49"),
   103 => (x"c0",x"f0",x"ea",x"87"),
   104 => (x"d0",x"87",x"c7",x"de"),
   105 => (x"49",x"c0",x"f0",x"e1"),
   106 => (x"87",x"c7",x"87",x"c8"),
   107 => (x"e7",x"49",x"c0",x"f0"),
   108 => (x"d8",x"87",x"73",x"49"),
   109 => (x"fb",x"f7",x"87",x"fe"),
   110 => (x"da",x"87",x"fb",x"ed"),
   111 => (x"87",x"38",x"33",x"32"),
   112 => (x"4f",x"53",x"44",x"41"),
   113 => (x"43",x"42",x"49",x"4e"),
   114 => (x"00",x"43",x"61",x"6e"),
   115 => (x"27",x"74",x"20",x"6c"),
   116 => (x"6f",x"61",x"64",x"20"),
   117 => (x"66",x"69",x"72",x"6d"),
   118 => (x"77",x"61",x"72",x"65"),
   119 => (x"0a",x"00",x"55",x"6e"),
   120 => (x"61",x"62",x"6c",x"65"),
   121 => (x"20",x"74",x"6f",x"20"),
   122 => (x"6c",x"6f",x"63",x"61"),
   123 => (x"74",x"65",x"20",x"70"),
   124 => (x"61",x"72",x"74",x"69"),
   125 => (x"74",x"69",x"6f",x"6e"),
   126 => (x"0a",x"00",x"48",x"75"),
   127 => (x"6e",x"74",x"69",x"6e"),
   128 => (x"67",x"20",x"66",x"6f"),
   129 => (x"72",x"20",x"70",x"61"),
   130 => (x"72",x"74",x"69",x"74"),
   131 => (x"69",x"6f",x"6e",x"0a"),
   132 => (x"00",x"49",x"6e",x"69"),
   133 => (x"74",x"69",x"61",x"6c"),
   134 => (x"69",x"7a",x"69",x"6e"),
   135 => (x"67",x"20",x"53",x"44"),
   136 => (x"20",x"63",x"61",x"72"),
   137 => (x"64",x"0a",x"00",x"46"),
   138 => (x"61",x"69",x"6c",x"65"),
   139 => (x"64",x"20",x"74",x"6f"),
   140 => (x"20",x"69",x"6e",x"69"),
   141 => (x"74",x"69",x"61",x"6c"),
   142 => (x"69",x"7a",x"65",x"20"),
   143 => (x"53",x"44",x"20",x"63"),
   144 => (x"61",x"72",x"64",x"0a"),
   145 => (x"00",x"00",x"00",x"00"),
   146 => (x"00",x"00",x"00",x"00"),
   147 => (x"08",x"33",x"fc",x"0f"),
   148 => (x"ff",x"00",x"df",x"f1"),
   149 => (x"80",x"60",x"f6",x"00"),
   150 => (x"00",x"00",x"12",x"1e"),
   151 => (x"e4",x"86",x"e3",x"48"),
   152 => (x"c3",x"ff",x"50",x"e3"),
   153 => (x"97",x"bf",x"48",x"c4"),
   154 => (x"a6",x"58",x"6e",x"49"),
   155 => (x"c3",x"ff",x"99",x"e3"),
   156 => (x"48",x"c3",x"ff",x"50"),
   157 => (x"c8",x"31",x"e3",x"97"),
   158 => (x"bf",x"48",x"c8",x"a6"),
   159 => (x"58",x"c4",x"66",x"48"),
   160 => (x"c3",x"ff",x"98",x"cc"),
   161 => (x"a6",x"58",x"c8",x"66"),
   162 => (x"b1",x"e3",x"48",x"c3"),
   163 => (x"ff",x"50",x"c8",x"31"),
   164 => (x"e3",x"97",x"bf",x"48"),
   165 => (x"d0",x"a6",x"58",x"cc"),
   166 => (x"66",x"48",x"c3",x"ff"),
   167 => (x"98",x"d4",x"a6",x"58"),
   168 => (x"d0",x"66",x"b1",x"e3"),
   169 => (x"48",x"c3",x"ff",x"50"),
   170 => (x"c8",x"31",x"e3",x"97"),
   171 => (x"bf",x"48",x"d8",x"a6"),
   172 => (x"58",x"d4",x"66",x"48"),
   173 => (x"c3",x"ff",x"98",x"dc"),
   174 => (x"a6",x"58",x"d8",x"66"),
   175 => (x"b1",x"71",x"48",x"e4"),
   176 => (x"8e",x"26",x"4f",x"0e"),
   177 => (x"5e",x"5b",x"5c",x"0e"),
   178 => (x"1e",x"71",x"4a",x"72"),
   179 => (x"49",x"c3",x"ff",x"99"),
   180 => (x"e3",x"09",x"97",x"79"),
   181 => (x"09",x"c1",x"c4",x"e0"),
   182 => (x"bf",x"05",x"c8",x"87"),
   183 => (x"d0",x"66",x"48",x"c9"),
   184 => (x"30",x"d4",x"a6",x"58"),
   185 => (x"d0",x"66",x"49",x"d8"),
   186 => (x"29",x"c3",x"ff",x"99"),
   187 => (x"e3",x"09",x"97",x"79"),
   188 => (x"09",x"d0",x"66",x"49"),
   189 => (x"d0",x"29",x"c3",x"ff"),
   190 => (x"99",x"e3",x"09",x"97"),
   191 => (x"79",x"09",x"d0",x"66"),
   192 => (x"49",x"c8",x"29",x"c3"),
   193 => (x"ff",x"99",x"e3",x"09"),
   194 => (x"97",x"79",x"09",x"d0"),
   195 => (x"66",x"49",x"c3",x"ff"),
   196 => (x"99",x"e3",x"09",x"97"),
   197 => (x"79",x"09",x"72",x"49"),
   198 => (x"d0",x"29",x"c3",x"ff"),
   199 => (x"99",x"e3",x"09",x"97"),
   200 => (x"79",x"09",x"97",x"bf"),
   201 => (x"48",x"c4",x"a6",x"58"),
   202 => (x"6e",x"4b",x"c3",x"ff"),
   203 => (x"9b",x"c9",x"f0",x"ff"),
   204 => (x"4c",x"c3",x"ff",x"ab"),
   205 => (x"05",x"dc",x"87",x"e3"),
   206 => (x"48",x"c3",x"ff",x"50"),
   207 => (x"e3",x"97",x"bf",x"48"),
   208 => (x"c4",x"a6",x"58",x"6e"),
   209 => (x"4b",x"c3",x"ff",x"9b"),
   210 => (x"c1",x"8c",x"02",x"c6"),
   211 => (x"87",x"c3",x"ff",x"ab"),
   212 => (x"02",x"e4",x"87",x"73"),
   213 => (x"4a",x"c4",x"b7",x"2a"),
   214 => (x"c0",x"f0",x"a2",x"49"),
   215 => (x"c0",x"e9",x"e0",x"87"),
   216 => (x"73",x"4a",x"cf",x"9a"),
   217 => (x"c0",x"f0",x"a2",x"49"),
   218 => (x"c0",x"e9",x"d4",x"87"),
   219 => (x"73",x"48",x"26",x"c2"),
   220 => (x"87",x"26",x"4d",x"26"),
   221 => (x"4c",x"26",x"4b",x"26"),
   222 => (x"4f",x"1e",x"c0",x"49"),
   223 => (x"e3",x"48",x"c3",x"ff"),
   224 => (x"50",x"c1",x"81",x"c3"),
   225 => (x"c8",x"b7",x"a9",x"04"),
   226 => (x"f2",x"87",x"26",x"4f"),
   227 => (x"1e",x"73",x"1e",x"e8"),
   228 => (x"87",x"c4",x"f8",x"df"),
   229 => (x"4b",x"c0",x"1e",x"c0"),
   230 => (x"ff",x"f0",x"c1",x"f7"),
   231 => (x"49",x"fc",x"e3",x"87"),
   232 => (x"c4",x"86",x"c1",x"a8"),
   233 => (x"05",x"c0",x"e8",x"87"),
   234 => (x"e3",x"48",x"c3",x"ff"),
   235 => (x"50",x"c1",x"c0",x"c0"),
   236 => (x"c0",x"c0",x"c0",x"1e"),
   237 => (x"c0",x"e1",x"f0",x"c1"),
   238 => (x"e9",x"49",x"fc",x"c6"),
   239 => (x"87",x"c4",x"86",x"70"),
   240 => (x"98",x"05",x"c9",x"87"),
   241 => (x"e3",x"48",x"c3",x"ff"),
   242 => (x"50",x"c1",x"48",x"cb"),
   243 => (x"87",x"fe",x"e9",x"87"),
   244 => (x"c1",x"8b",x"05",x"fe"),
   245 => (x"ff",x"87",x"c0",x"48"),
   246 => (x"fe",x"da",x"87",x"43"),
   247 => (x"4d",x"44",x"34",x"31"),
   248 => (x"20",x"25",x"64",x"0a"),
   249 => (x"00",x"43",x"4d",x"44"),
   250 => (x"35",x"35",x"20",x"25"),
   251 => (x"64",x"0a",x"00",x"43"),
   252 => (x"4d",x"44",x"34",x"31"),
   253 => (x"20",x"25",x"64",x"0a"),
   254 => (x"00",x"43",x"4d",x"44"),
   255 => (x"35",x"35",x"20",x"25"),
   256 => (x"64",x"0a",x"00",x"69"),
   257 => (x"6e",x"69",x"74",x"20"),
   258 => (x"25",x"64",x"0a",x"20"),
   259 => (x"20",x"00",x"69",x"6e"),
   260 => (x"69",x"74",x"20",x"25"),
   261 => (x"64",x"0a",x"20",x"20"),
   262 => (x"00",x"43",x"6d",x"64"),
   263 => (x"5f",x"69",x"6e",x"69"),
   264 => (x"74",x"0a",x"00",x"43"),
   265 => (x"4d",x"44",x"38",x"5f"),
   266 => (x"34",x"20",x"72",x"65"),
   267 => (x"73",x"70",x"6f",x"6e"),
   268 => (x"73",x"65",x"3a",x"20"),
   269 => (x"25",x"64",x"0a",x"00"),
   270 => (x"43",x"4d",x"44",x"35"),
   271 => (x"38",x"20",x"25",x"64"),
   272 => (x"0a",x"20",x"20",x"00"),
   273 => (x"43",x"4d",x"44",x"35"),
   274 => (x"38",x"5f",x"32",x"20"),
   275 => (x"25",x"64",x"0a",x"20"),
   276 => (x"20",x"00",x"43",x"4d"),
   277 => (x"44",x"35",x"38",x"20"),
   278 => (x"25",x"64",x"0a",x"20"),
   279 => (x"20",x"00",x"53",x"44"),
   280 => (x"48",x"43",x"20",x"49"),
   281 => (x"6e",x"69",x"74",x"69"),
   282 => (x"61",x"6c",x"69",x"7a"),
   283 => (x"61",x"74",x"69",x"6f"),
   284 => (x"6e",x"20",x"65",x"72"),
   285 => (x"72",x"6f",x"72",x"21"),
   286 => (x"0a",x"00",x"63",x"6d"),
   287 => (x"64",x"5f",x"43",x"4d"),
   288 => (x"44",x"38",x"20",x"72"),
   289 => (x"65",x"73",x"70",x"6f"),
   290 => (x"6e",x"73",x"65",x"3a"),
   291 => (x"20",x"25",x"64",x"0a"),
   292 => (x"00",x"52",x"65",x"61"),
   293 => (x"64",x"20",x"63",x"6f"),
   294 => (x"6d",x"6d",x"61",x"6e"),
   295 => (x"64",x"20",x"66",x"61"),
   296 => (x"69",x"6c",x"65",x"64"),
   297 => (x"20",x"61",x"74",x"20"),
   298 => (x"25",x"64",x"20",x"28"),
   299 => (x"25",x"64",x"29",x"0a"),
   300 => (x"00",x"1e",x"73",x"1e"),
   301 => (x"e3",x"48",x"c3",x"ff"),
   302 => (x"50",x"d0",x"d9",x"49"),
   303 => (x"c0",x"e4",x"ca",x"87"),
   304 => (x"d3",x"4b",x"c0",x"1e"),
   305 => (x"c0",x"ff",x"f0",x"c1"),
   306 => (x"c1",x"49",x"f7",x"f6"),
   307 => (x"87",x"c4",x"86",x"70"),
   308 => (x"98",x"05",x"c9",x"87"),
   309 => (x"e3",x"48",x"c3",x"ff"),
   310 => (x"50",x"c1",x"48",x"cb"),
   311 => (x"87",x"fa",x"d9",x"87"),
   312 => (x"c1",x"8b",x"05",x"ff"),
   313 => (x"dc",x"87",x"c0",x"48"),
   314 => (x"fa",x"ca",x"87",x"1e"),
   315 => (x"73",x"1e",x"1e",x"fa"),
   316 => (x"c7",x"87",x"c6",x"ea"),
   317 => (x"1e",x"c0",x"e1",x"f0"),
   318 => (x"c1",x"c8",x"49",x"f7"),
   319 => (x"c5",x"87",x"70",x"4b"),
   320 => (x"73",x"1e",x"d1",x"fa"),
   321 => (x"1e",x"c0",x"ee",x"de"),
   322 => (x"87",x"cc",x"86",x"c1"),
   323 => (x"ab",x"02",x"c8",x"87"),
   324 => (x"fe",x"de",x"87",x"c0"),
   325 => (x"48",x"c1",x"ff",x"87"),
   326 => (x"f5",x"c0",x"87",x"70"),
   327 => (x"49",x"cf",x"ff",x"ff"),
   328 => (x"99",x"c6",x"ea",x"a9"),
   329 => (x"02",x"c8",x"87",x"fe"),
   330 => (x"c7",x"87",x"c0",x"48"),
   331 => (x"c1",x"e8",x"87",x"e3"),
   332 => (x"48",x"c3",x"ff",x"50"),
   333 => (x"c0",x"f1",x"4b",x"f9"),
   334 => (x"d2",x"87",x"70",x"98"),
   335 => (x"02",x"c1",x"c6",x"87"),
   336 => (x"c0",x"1e",x"c0",x"ff"),
   337 => (x"f0",x"c1",x"fa",x"49"),
   338 => (x"f5",x"f8",x"87",x"c4"),
   339 => (x"86",x"70",x"98",x"05"),
   340 => (x"c0",x"f3",x"87",x"e3"),
   341 => (x"48",x"c3",x"ff",x"50"),
   342 => (x"e3",x"97",x"bf",x"48"),
   343 => (x"c4",x"a6",x"58",x"6e"),
   344 => (x"49",x"c3",x"ff",x"99"),
   345 => (x"e3",x"48",x"c3",x"ff"),
   346 => (x"50",x"e3",x"48",x"c3"),
   347 => (x"ff",x"50",x"e3",x"48"),
   348 => (x"c3",x"ff",x"50",x"e3"),
   349 => (x"48",x"c3",x"ff",x"50"),
   350 => (x"c1",x"c0",x"99",x"02"),
   351 => (x"c4",x"87",x"c1",x"48"),
   352 => (x"d5",x"87",x"c0",x"48"),
   353 => (x"d1",x"87",x"c2",x"ab"),
   354 => (x"05",x"c4",x"87",x"c0"),
   355 => (x"48",x"c8",x"87",x"c1"),
   356 => (x"8b",x"05",x"fe",x"e2"),
   357 => (x"87",x"c0",x"48",x"26"),
   358 => (x"f7",x"da",x"87",x"1e"),
   359 => (x"73",x"1e",x"c1",x"c4"),
   360 => (x"e0",x"48",x"c1",x"78"),
   361 => (x"eb",x"48",x"c3",x"ef"),
   362 => (x"50",x"c7",x"4b",x"e7"),
   363 => (x"48",x"c3",x"50",x"f7"),
   364 => (x"c7",x"87",x"e7",x"48"),
   365 => (x"c2",x"50",x"e3",x"48"),
   366 => (x"c3",x"ff",x"50",x"c0"),
   367 => (x"1e",x"c0",x"e5",x"d0"),
   368 => (x"c1",x"c0",x"49",x"f3"),
   369 => (x"fd",x"87",x"c4",x"86"),
   370 => (x"c1",x"a8",x"05",x"c2"),
   371 => (x"87",x"c1",x"4b",x"c2"),
   372 => (x"ab",x"05",x"c5",x"87"),
   373 => (x"c0",x"48",x"c0",x"f1"),
   374 => (x"87",x"c1",x"8b",x"05"),
   375 => (x"ff",x"cc",x"87",x"fc"),
   376 => (x"c9",x"87",x"c1",x"c4"),
   377 => (x"e4",x"58",x"c1",x"c4"),
   378 => (x"e0",x"bf",x"05",x"cd"),
   379 => (x"87",x"c1",x"1e",x"c0"),
   380 => (x"ff",x"f0",x"c1",x"d0"),
   381 => (x"49",x"f3",x"cb",x"87"),
   382 => (x"c4",x"86",x"e3",x"48"),
   383 => (x"c3",x"ff",x"50",x"e7"),
   384 => (x"48",x"c3",x"50",x"e3"),
   385 => (x"48",x"c3",x"ff",x"50"),
   386 => (x"c1",x"48",x"f5",x"e8"),
   387 => (x"87",x"0e",x"5e",x"5b"),
   388 => (x"5c",x"5d",x"0e",x"1e"),
   389 => (x"71",x"4a",x"c0",x"4d"),
   390 => (x"e3",x"48",x"c3",x"ff"),
   391 => (x"50",x"e7",x"48",x"c2"),
   392 => (x"50",x"eb",x"48",x"c7"),
   393 => (x"50",x"e3",x"48",x"c3"),
   394 => (x"ff",x"50",x"72",x"1e"),
   395 => (x"c0",x"ff",x"f0",x"c1"),
   396 => (x"d1",x"49",x"f2",x"ce"),
   397 => (x"87",x"c4",x"86",x"70"),
   398 => (x"98",x"05",x"c1",x"c9"),
   399 => (x"87",x"c5",x"ee",x"cd"),
   400 => (x"df",x"4b",x"e3",x"48"),
   401 => (x"c3",x"ff",x"50",x"e3"),
   402 => (x"97",x"bf",x"48",x"c4"),
   403 => (x"a6",x"58",x"6e",x"49"),
   404 => (x"c3",x"ff",x"99",x"c3"),
   405 => (x"fe",x"a9",x"05",x"de"),
   406 => (x"87",x"c0",x"4c",x"ef"),
   407 => (x"fd",x"87",x"d4",x"66"),
   408 => (x"08",x"78",x"08",x"d4"),
   409 => (x"66",x"48",x"c4",x"80"),
   410 => (x"d8",x"a6",x"58",x"c1"),
   411 => (x"84",x"c2",x"c0",x"b7"),
   412 => (x"ac",x"04",x"e7",x"87"),
   413 => (x"c1",x"4b",x"4d",x"c1"),
   414 => (x"8b",x"05",x"ff",x"c5"),
   415 => (x"87",x"e3",x"48",x"c3"),
   416 => (x"ff",x"50",x"e7",x"48"),
   417 => (x"c3",x"50",x"75",x"48"),
   418 => (x"26",x"f3",x"e5",x"87"),
   419 => (x"1e",x"73",x"1e",x"71"),
   420 => (x"4b",x"73",x"49",x"d8"),
   421 => (x"29",x"c3",x"ff",x"99"),
   422 => (x"73",x"4a",x"c8",x"2a"),
   423 => (x"cf",x"fc",x"c0",x"9a"),
   424 => (x"72",x"b1",x"73",x"4a"),
   425 => (x"c8",x"32",x"c0",x"ff"),
   426 => (x"f0",x"c0",x"c0",x"9a"),
   427 => (x"72",x"b1",x"73",x"4a"),
   428 => (x"d8",x"32",x"ff",x"c0"),
   429 => (x"c0",x"c0",x"c0",x"9a"),
   430 => (x"72",x"b1",x"71",x"48"),
   431 => (x"c4",x"87",x"26",x"4d"),
   432 => (x"26",x"4c",x"26",x"4b"),
   433 => (x"26",x"4f",x"1e",x"73"),
   434 => (x"1e",x"71",x"4b",x"73"),
   435 => (x"49",x"c8",x"29",x"c3"),
   436 => (x"ff",x"99",x"73",x"4a"),
   437 => (x"c8",x"32",x"cf",x"fc"),
   438 => (x"c0",x"9a",x"72",x"b1"),
   439 => (x"71",x"48",x"e2",x"87"),
   440 => (x"0e",x"5e",x"5b",x"5c"),
   441 => (x"0e",x"71",x"4b",x"c0"),
   442 => (x"4c",x"d0",x"66",x"48"),
   443 => (x"c0",x"b7",x"a8",x"06"),
   444 => (x"c0",x"e3",x"87",x"13"),
   445 => (x"4a",x"cc",x"66",x"97"),
   446 => (x"bf",x"49",x"cc",x"66"),
   447 => (x"48",x"c1",x"80",x"d0"),
   448 => (x"a6",x"58",x"71",x"b7"),
   449 => (x"aa",x"02",x"c4",x"87"),
   450 => (x"c1",x"48",x"cc",x"87"),
   451 => (x"c1",x"84",x"d0",x"66"),
   452 => (x"b7",x"ac",x"04",x"ff"),
   453 => (x"dd",x"87",x"c0",x"48"),
   454 => (x"c2",x"87",x"26",x"4d"),
   455 => (x"26",x"4c",x"26",x"4b"),
   456 => (x"26",x"4f",x"0e",x"5e"),
   457 => (x"5b",x"5c",x"0e",x"1e"),
   458 => (x"c1",x"cd",x"e2",x"48"),
   459 => (x"ff",x"78",x"c1",x"cc"),
   460 => (x"f2",x"48",x"c0",x"78"),
   461 => (x"c0",x"ea",x"c7",x"49"),
   462 => (x"da",x"cf",x"87",x"c1"),
   463 => (x"c4",x"ea",x"1e",x"c0"),
   464 => (x"49",x"fb",x"c9",x"87"),
   465 => (x"c4",x"86",x"70",x"98"),
   466 => (x"05",x"c5",x"87",x"c0"),
   467 => (x"48",x"ca",x"f0",x"87"),
   468 => (x"c0",x"4b",x"c1",x"cd"),
   469 => (x"de",x"48",x"c1",x"78"),
   470 => (x"c8",x"1e",x"c0",x"ea"),
   471 => (x"d4",x"1e",x"c1",x"c5"),
   472 => (x"e0",x"49",x"fd",x"fb"),
   473 => (x"87",x"c8",x"86",x"70"),
   474 => (x"98",x"05",x"c6",x"87"),
   475 => (x"c1",x"cd",x"de",x"48"),
   476 => (x"c0",x"78",x"c8",x"1e"),
   477 => (x"c0",x"ea",x"dd",x"1e"),
   478 => (x"c1",x"c5",x"fc",x"49"),
   479 => (x"fd",x"e1",x"87",x"c8"),
   480 => (x"86",x"70",x"98",x"05"),
   481 => (x"c6",x"87",x"c1",x"cd"),
   482 => (x"de",x"48",x"c0",x"78"),
   483 => (x"c8",x"1e",x"c0",x"ea"),
   484 => (x"e6",x"1e",x"c1",x"c5"),
   485 => (x"fc",x"49",x"fd",x"c7"),
   486 => (x"87",x"c8",x"86",x"70"),
   487 => (x"98",x"05",x"c5",x"87"),
   488 => (x"c0",x"48",x"c9",x"db"),
   489 => (x"87",x"c1",x"cd",x"de"),
   490 => (x"bf",x"1e",x"c0",x"ea"),
   491 => (x"ef",x"1e",x"c0",x"e3"),
   492 => (x"f5",x"87",x"c8",x"86"),
   493 => (x"c1",x"cd",x"de",x"bf"),
   494 => (x"02",x"c1",x"ed",x"87"),
   495 => (x"c1",x"c4",x"ea",x"4a"),
   496 => (x"48",x"c6",x"fe",x"a0"),
   497 => (x"4c",x"c1",x"cb",x"f0"),
   498 => (x"bf",x"4b",x"c1",x"cc"),
   499 => (x"e8",x"9f",x"bf",x"49"),
   500 => (x"c4",x"a6",x"5a",x"c5"),
   501 => (x"d6",x"ea",x"a9",x"05"),
   502 => (x"c0",x"cc",x"87",x"c8"),
   503 => (x"a4",x"4a",x"6a",x"49"),
   504 => (x"fa",x"e9",x"87",x"70"),
   505 => (x"4b",x"db",x"87",x"c7"),
   506 => (x"fe",x"a2",x"49",x"9f"),
   507 => (x"69",x"49",x"ca",x"e9"),
   508 => (x"d5",x"a9",x"02",x"c0"),
   509 => (x"cc",x"87",x"c0",x"e8"),
   510 => (x"c4",x"49",x"d7",x"cd"),
   511 => (x"87",x"c0",x"48",x"c7"),
   512 => (x"fe",x"87",x"73",x"1e"),
   513 => (x"c0",x"e8",x"e2",x"1e"),
   514 => (x"c0",x"e2",x"db",x"87"),
   515 => (x"c1",x"c4",x"ea",x"1e"),
   516 => (x"73",x"49",x"f7",x"f8"),
   517 => (x"87",x"cc",x"86",x"70"),
   518 => (x"98",x"05",x"c0",x"c5"),
   519 => (x"87",x"c0",x"48",x"c7"),
   520 => (x"de",x"87",x"c0",x"e8"),
   521 => (x"fa",x"49",x"d6",x"e1"),
   522 => (x"87",x"c0",x"eb",x"c2"),
   523 => (x"1e",x"c0",x"e1",x"f6"),
   524 => (x"87",x"c8",x"1e",x"c0"),
   525 => (x"eb",x"da",x"1e",x"c1"),
   526 => (x"c5",x"fc",x"49",x"fa"),
   527 => (x"e2",x"87",x"cc",x"86"),
   528 => (x"70",x"98",x"05",x"c0"),
   529 => (x"c9",x"87",x"c1",x"cc"),
   530 => (x"f2",x"48",x"c1",x"78"),
   531 => (x"c0",x"e4",x"87",x"c8"),
   532 => (x"1e",x"c0",x"eb",x"e3"),
   533 => (x"1e",x"c1",x"c5",x"e0"),
   534 => (x"49",x"fa",x"c4",x"87"),
   535 => (x"c8",x"86",x"70",x"98"),
   536 => (x"02",x"c0",x"cf",x"87"),
   537 => (x"c0",x"e9",x"e1",x"1e"),
   538 => (x"c0",x"e0",x"fb",x"87"),
   539 => (x"c4",x"86",x"c0",x"48"),
   540 => (x"c6",x"cd",x"87",x"c1"),
   541 => (x"cc",x"e8",x"97",x"bf"),
   542 => (x"49",x"c1",x"d5",x"a9"),
   543 => (x"05",x"c0",x"cd",x"87"),
   544 => (x"c1",x"cc",x"e9",x"97"),
   545 => (x"bf",x"49",x"c2",x"ea"),
   546 => (x"a9",x"02",x"c0",x"c5"),
   547 => (x"87",x"c0",x"48",x"c5"),
   548 => (x"ee",x"87",x"c1",x"c4"),
   549 => (x"ea",x"97",x"bf",x"49"),
   550 => (x"c3",x"e9",x"a9",x"02"),
   551 => (x"c0",x"d2",x"87",x"c1"),
   552 => (x"c4",x"ea",x"97",x"bf"),
   553 => (x"49",x"c3",x"eb",x"a9"),
   554 => (x"02",x"c0",x"c5",x"87"),
   555 => (x"c0",x"48",x"c5",x"cf"),
   556 => (x"87",x"c1",x"c4",x"f5"),
   557 => (x"97",x"bf",x"49",x"71"),
   558 => (x"99",x"05",x"c0",x"cc"),
   559 => (x"87",x"c1",x"c4",x"f6"),
   560 => (x"97",x"bf",x"49",x"c2"),
   561 => (x"a9",x"02",x"c0",x"c5"),
   562 => (x"87",x"c0",x"48",x"c4"),
   563 => (x"f2",x"87",x"c1",x"c4"),
   564 => (x"f7",x"97",x"bf",x"48"),
   565 => (x"c1",x"cc",x"ee",x"58"),
   566 => (x"c1",x"cc",x"ea",x"bf"),
   567 => (x"48",x"c1",x"88",x"c1"),
   568 => (x"cc",x"f2",x"58",x"c1"),
   569 => (x"c4",x"f8",x"97",x"bf"),
   570 => (x"49",x"73",x"81",x"c1"),
   571 => (x"c4",x"f9",x"97",x"bf"),
   572 => (x"4a",x"c8",x"32",x"c1"),
   573 => (x"cc",x"fe",x"48",x"72"),
   574 => (x"a1",x"78",x"c1",x"c4"),
   575 => (x"fa",x"97",x"bf",x"48"),
   576 => (x"c1",x"cd",x"d6",x"58"),
   577 => (x"c1",x"cc",x"f2",x"bf"),
   578 => (x"02",x"c2",x"e2",x"87"),
   579 => (x"c8",x"1e",x"c0",x"e9"),
   580 => (x"fe",x"1e",x"c1",x"c5"),
   581 => (x"fc",x"49",x"f7",x"c7"),
   582 => (x"87",x"c8",x"86",x"70"),
   583 => (x"98",x"02",x"c0",x"c5"),
   584 => (x"87",x"c0",x"48",x"c3"),
   585 => (x"da",x"87",x"c1",x"cc"),
   586 => (x"ea",x"bf",x"48",x"c4"),
   587 => (x"30",x"c1",x"cd",x"da"),
   588 => (x"58",x"c1",x"cc",x"ea"),
   589 => (x"bf",x"4a",x"c1",x"cd"),
   590 => (x"d2",x"5a",x"c1",x"c5"),
   591 => (x"cf",x"97",x"bf",x"49"),
   592 => (x"c8",x"31",x"c1",x"c5"),
   593 => (x"ce",x"97",x"bf",x"4b"),
   594 => (x"73",x"a1",x"49",x"c1"),
   595 => (x"c5",x"d0",x"97",x"bf"),
   596 => (x"4b",x"d0",x"33",x"73"),
   597 => (x"a1",x"49",x"c1",x"c5"),
   598 => (x"d1",x"97",x"bf",x"4b"),
   599 => (x"d8",x"33",x"73",x"a1"),
   600 => (x"49",x"c1",x"cd",x"de"),
   601 => (x"59",x"c1",x"cd",x"d2"),
   602 => (x"bf",x"91",x"c1",x"cc"),
   603 => (x"fe",x"bf",x"81",x"c1"),
   604 => (x"cd",x"c6",x"59",x"c1"),
   605 => (x"c5",x"d7",x"97",x"bf"),
   606 => (x"4b",x"c8",x"33",x"c1"),
   607 => (x"c5",x"d6",x"97",x"bf"),
   608 => (x"4c",x"74",x"a3",x"4b"),
   609 => (x"c1",x"c5",x"d8",x"97"),
   610 => (x"bf",x"4c",x"d0",x"34"),
   611 => (x"74",x"a3",x"4b",x"c1"),
   612 => (x"c5",x"d9",x"97",x"bf"),
   613 => (x"4c",x"cf",x"9c",x"d8"),
   614 => (x"34",x"74",x"a3",x"4b"),
   615 => (x"c1",x"cd",x"ca",x"5b"),
   616 => (x"c2",x"8b",x"73",x"92"),
   617 => (x"c1",x"cd",x"ca",x"48"),
   618 => (x"72",x"a1",x"78",x"c1"),
   619 => (x"d0",x"87",x"c1",x"c4"),
   620 => (x"fc",x"97",x"bf",x"49"),
   621 => (x"c8",x"31",x"c1",x"c4"),
   622 => (x"fb",x"97",x"bf",x"4a"),
   623 => (x"72",x"a1",x"49",x"c1"),
   624 => (x"cd",x"da",x"59",x"c5"),
   625 => (x"31",x"c7",x"ff",x"81"),
   626 => (x"c9",x"29",x"c1",x"cd"),
   627 => (x"d2",x"59",x"c1",x"c5"),
   628 => (x"c1",x"97",x"bf",x"4a"),
   629 => (x"c8",x"32",x"c1",x"c5"),
   630 => (x"c0",x"97",x"bf",x"4b"),
   631 => (x"73",x"a2",x"4a",x"c1"),
   632 => (x"cd",x"de",x"5a",x"c1"),
   633 => (x"cd",x"d2",x"bf",x"92"),
   634 => (x"c1",x"cc",x"fe",x"bf"),
   635 => (x"82",x"c1",x"cd",x"ce"),
   636 => (x"5a",x"c1",x"cd",x"c6"),
   637 => (x"48",x"c0",x"78",x"c1"),
   638 => (x"cd",x"c2",x"48",x"72"),
   639 => (x"a1",x"78",x"c1",x"48"),
   640 => (x"26",x"f4",x"d8",x"87"),
   641 => (x"4e",x"6f",x"20",x"70"),
   642 => (x"61",x"72",x"74",x"69"),
   643 => (x"74",x"69",x"6f",x"6e"),
   644 => (x"20",x"73",x"69",x"67"),
   645 => (x"6e",x"61",x"74",x"75"),
   646 => (x"72",x"65",x"20",x"66"),
   647 => (x"6f",x"75",x"6e",x"64"),
   648 => (x"0a",x"00",x"52",x"65"),
   649 => (x"61",x"64",x"69",x"6e"),
   650 => (x"67",x"20",x"62",x"6f"),
   651 => (x"6f",x"74",x"20",x"73"),
   652 => (x"65",x"63",x"74",x"6f"),
   653 => (x"72",x"20",x"25",x"64"),
   654 => (x"0a",x"00",x"52",x"65"),
   655 => (x"61",x"64",x"20",x"62"),
   656 => (x"6f",x"6f",x"74",x"20"),
   657 => (x"73",x"65",x"63",x"74"),
   658 => (x"6f",x"72",x"20",x"66"),
   659 => (x"72",x"6f",x"6d",x"20"),
   660 => (x"66",x"69",x"72",x"73"),
   661 => (x"74",x"20",x"70",x"61"),
   662 => (x"72",x"74",x"69",x"74"),
   663 => (x"69",x"6f",x"6e",x"0a"),
   664 => (x"00",x"55",x"6e",x"73"),
   665 => (x"75",x"70",x"70",x"6f"),
   666 => (x"72",x"74",x"65",x"64"),
   667 => (x"20",x"70",x"61",x"72"),
   668 => (x"74",x"69",x"74",x"69"),
   669 => (x"6f",x"6e",x"20",x"74"),
   670 => (x"79",x"70",x"65",x"21"),
   671 => (x"0d",x"00",x"46",x"41"),
   672 => (x"54",x"33",x"32",x"20"),
   673 => (x"20",x"20",x"00",x"52"),
   674 => (x"65",x"61",x"64",x"69"),
   675 => (x"6e",x"67",x"20",x"4d"),
   676 => (x"42",x"52",x"0a",x"00"),
   677 => (x"46",x"41",x"54",x"31"),
   678 => (x"36",x"20",x"20",x"20"),
   679 => (x"00",x"46",x"41",x"54"),
   680 => (x"33",x"32",x"20",x"20"),
   681 => (x"20",x"00",x"46",x"41"),
   682 => (x"54",x"31",x"32",x"20"),
   683 => (x"20",x"20",x"00",x"50"),
   684 => (x"61",x"72",x"74",x"69"),
   685 => (x"74",x"69",x"6f",x"6e"),
   686 => (x"63",x"6f",x"75",x"6e"),
   687 => (x"74",x"20",x"25",x"64"),
   688 => (x"0a",x"00",x"48",x"75"),
   689 => (x"6e",x"74",x"69",x"6e"),
   690 => (x"67",x"20",x"66",x"6f"),
   691 => (x"72",x"20",x"66",x"69"),
   692 => (x"6c",x"65",x"73",x"79"),
   693 => (x"73",x"74",x"65",x"6d"),
   694 => (x"0a",x"00",x"46",x"41"),
   695 => (x"54",x"33",x"32",x"20"),
   696 => (x"20",x"20",x"00",x"46"),
   697 => (x"41",x"54",x"31",x"36"),
   698 => (x"20",x"20",x"20",x"00"),
   699 => (x"52",x"65",x"61",x"64"),
   700 => (x"69",x"6e",x"67",x"20"),
   701 => (x"64",x"69",x"72",x"65"),
   702 => (x"63",x"74",x"6f",x"72"),
   703 => (x"79",x"20",x"73",x"65"),
   704 => (x"63",x"74",x"6f",x"72"),
   705 => (x"20",x"25",x"64",x"0a"),
   706 => (x"00",x"66",x"69",x"6c"),
   707 => (x"65",x"20",x"22",x"25"),
   708 => (x"73",x"22",x"20",x"66"),
   709 => (x"6f",x"75",x"6e",x"64"),
   710 => (x"0d",x"00",x"47",x"65"),
   711 => (x"74",x"46",x"41",x"54"),
   712 => (x"4c",x"69",x"6e",x"6b"),
   713 => (x"20",x"72",x"65",x"74"),
   714 => (x"75",x"72",x"6e",x"65"),
   715 => (x"64",x"20",x"25",x"64"),
   716 => (x"0a",x"00",x"43",x"61"),
   717 => (x"6e",x"27",x"74",x"20"),
   718 => (x"6f",x"70",x"65",x"6e"),
   719 => (x"20",x"25",x"73",x"0a"),
   720 => (x"00",x"0e",x"5e",x"5b"),
   721 => (x"5c",x"5d",x"0e",x"71"),
   722 => (x"4a",x"c1",x"cc",x"f2"),
   723 => (x"bf",x"02",x"cc",x"87"),
   724 => (x"72",x"4b",x"c7",x"b7"),
   725 => (x"2b",x"72",x"4c",x"c1"),
   726 => (x"ff",x"9c",x"ca",x"87"),
   727 => (x"72",x"4b",x"c8",x"b7"),
   728 => (x"2b",x"72",x"4c",x"c3"),
   729 => (x"ff",x"9c",x"c1",x"cd"),
   730 => (x"e2",x"bf",x"ab",x"02"),
   731 => (x"de",x"87",x"c1",x"c4"),
   732 => (x"ea",x"1e",x"c1",x"cc"),
   733 => (x"fe",x"bf",x"49",x"73"),
   734 => (x"81",x"ea",x"d1",x"87"),
   735 => (x"c4",x"86",x"70",x"98"),
   736 => (x"05",x"c5",x"87",x"c0"),
   737 => (x"48",x"c0",x"f6",x"87"),
   738 => (x"c1",x"cd",x"e6",x"5b"),
   739 => (x"c1",x"cc",x"f2",x"bf"),
   740 => (x"02",x"d9",x"87",x"74"),
   741 => (x"4a",x"c4",x"92",x"c1"),
   742 => (x"c4",x"ea",x"82",x"6a"),
   743 => (x"49",x"eb",x"ec",x"87"),
   744 => (x"70",x"49",x"71",x"4d"),
   745 => (x"cf",x"ff",x"ff",x"ff"),
   746 => (x"ff",x"9d",x"d0",x"87"),
   747 => (x"74",x"4a",x"c2",x"92"),
   748 => (x"c1",x"c4",x"ea",x"82"),
   749 => (x"9f",x"6a",x"49",x"ec"),
   750 => (x"cc",x"87",x"70",x"4d"),
   751 => (x"75",x"48",x"ed",x"d9"),
   752 => (x"87",x"0e",x"5e",x"5b"),
   753 => (x"5c",x"5d",x"0e",x"f4"),
   754 => (x"86",x"71",x"4c",x"c0"),
   755 => (x"4b",x"c1",x"cd",x"e2"),
   756 => (x"48",x"ff",x"78",x"c1"),
   757 => (x"cd",x"c6",x"bf",x"4d"),
   758 => (x"c1",x"cd",x"ca",x"bf"),
   759 => (x"7e",x"c1",x"cc",x"f2"),
   760 => (x"bf",x"02",x"c9",x"87"),
   761 => (x"c1",x"cc",x"ea",x"bf"),
   762 => (x"4a",x"c4",x"32",x"c7"),
   763 => (x"87",x"c1",x"cd",x"ce"),
   764 => (x"bf",x"4a",x"c4",x"32"),
   765 => (x"c8",x"a6",x"5a",x"c8"),
   766 => (x"a6",x"48",x"c0",x"78"),
   767 => (x"c4",x"66",x"48",x"c0"),
   768 => (x"a8",x"06",x"c3",x"cf"),
   769 => (x"87",x"c8",x"66",x"49"),
   770 => (x"cf",x"99",x"05",x"c0"),
   771 => (x"e3",x"87",x"6e",x"1e"),
   772 => (x"c0",x"eb",x"ec",x"1e"),
   773 => (x"d2",x"d0",x"87",x"c1"),
   774 => (x"c4",x"ea",x"1e",x"cc"),
   775 => (x"66",x"49",x"48",x"c1"),
   776 => (x"80",x"d0",x"a6",x"58"),
   777 => (x"71",x"49",x"e7",x"e4"),
   778 => (x"87",x"cc",x"86",x"c1"),
   779 => (x"c4",x"ea",x"4b",x"c3"),
   780 => (x"87",x"c0",x"e0",x"83"),
   781 => (x"97",x"6b",x"49",x"71"),
   782 => (x"99",x"02",x"c2",x"c5"),
   783 => (x"87",x"97",x"6b",x"49"),
   784 => (x"c3",x"e5",x"a9",x"02"),
   785 => (x"c1",x"fb",x"87",x"cb"),
   786 => (x"a3",x"49",x"97",x"69"),
   787 => (x"49",x"d8",x"99",x"05"),
   788 => (x"c1",x"ef",x"87",x"cb"),
   789 => (x"1e",x"c0",x"e0",x"66"),
   790 => (x"1e",x"73",x"49",x"ea"),
   791 => (x"c2",x"87",x"c8",x"86"),
   792 => (x"70",x"98",x"05",x"c1"),
   793 => (x"dc",x"87",x"dc",x"a3"),
   794 => (x"4a",x"6a",x"49",x"e8"),
   795 => (x"de",x"87",x"70",x"4a"),
   796 => (x"c4",x"a4",x"49",x"72"),
   797 => (x"79",x"da",x"a3",x"4a"),
   798 => (x"9f",x"6a",x"49",x"e9"),
   799 => (x"c8",x"87",x"c4",x"a6"),
   800 => (x"58",x"c1",x"cc",x"f2"),
   801 => (x"bf",x"02",x"d8",x"87"),
   802 => (x"d4",x"a3",x"4a",x"9f"),
   803 => (x"6a",x"49",x"e8",x"f5"),
   804 => (x"87",x"70",x"49",x"c0"),
   805 => (x"ff",x"ff",x"99",x"71"),
   806 => (x"48",x"d0",x"30",x"c8"),
   807 => (x"a6",x"58",x"c5",x"87"),
   808 => (x"c4",x"a6",x"48",x"c0"),
   809 => (x"78",x"c4",x"66",x"4a"),
   810 => (x"6e",x"82",x"c8",x"a4"),
   811 => (x"49",x"72",x"79",x"c0"),
   812 => (x"7c",x"dc",x"66",x"1e"),
   813 => (x"c0",x"ec",x"c9",x"1e"),
   814 => (x"cf",x"ec",x"87",x"c8"),
   815 => (x"86",x"c1",x"48",x"c1"),
   816 => (x"d0",x"87",x"c8",x"66"),
   817 => (x"48",x"c1",x"80",x"cc"),
   818 => (x"a6",x"58",x"c8",x"66"),
   819 => (x"48",x"c4",x"66",x"a8"),
   820 => (x"04",x"fc",x"f1",x"87"),
   821 => (x"c1",x"cc",x"f2",x"bf"),
   822 => (x"02",x"c0",x"f4",x"87"),
   823 => (x"75",x"49",x"f9",x"e0"),
   824 => (x"87",x"70",x"4d",x"75"),
   825 => (x"1e",x"c0",x"ec",x"da"),
   826 => (x"1e",x"ce",x"fb",x"87"),
   827 => (x"c8",x"86",x"75",x"49"),
   828 => (x"cf",x"ff",x"ff",x"ff"),
   829 => (x"f8",x"99",x"a9",x"02"),
   830 => (x"d6",x"87",x"75",x"49"),
   831 => (x"c2",x"89",x"c1",x"cc"),
   832 => (x"ea",x"bf",x"91",x"c1"),
   833 => (x"cd",x"c2",x"bf",x"48"),
   834 => (x"71",x"80",x"c4",x"a6"),
   835 => (x"58",x"fb",x"e7",x"87"),
   836 => (x"c0",x"48",x"f4",x"8e"),
   837 => (x"e8",x"c3",x"87",x"0e"),
   838 => (x"5e",x"5b",x"5c",x"5d"),
   839 => (x"0e",x"1e",x"71",x"4b"),
   840 => (x"73",x"1e",x"c1",x"cd"),
   841 => (x"e6",x"49",x"fa",x"d8"),
   842 => (x"87",x"c4",x"86",x"70"),
   843 => (x"98",x"02",x"c1",x"f7"),
   844 => (x"87",x"c1",x"cd",x"ea"),
   845 => (x"bf",x"49",x"c7",x"ff"),
   846 => (x"81",x"c9",x"29",x"c4"),
   847 => (x"a6",x"59",x"c0",x"4d"),
   848 => (x"4c",x"6e",x"48",x"c0"),
   849 => (x"b7",x"a8",x"06",x"c1"),
   850 => (x"ed",x"87",x"c1",x"cd"),
   851 => (x"c2",x"bf",x"49",x"c1"),
   852 => (x"cd",x"ee",x"bf",x"4a"),
   853 => (x"c2",x"8a",x"c1",x"cc"),
   854 => (x"ea",x"bf",x"92",x"72"),
   855 => (x"a1",x"49",x"c1",x"cc"),
   856 => (x"ee",x"bf",x"4a",x"74"),
   857 => (x"9a",x"72",x"a1",x"49"),
   858 => (x"d4",x"66",x"1e",x"71"),
   859 => (x"49",x"e2",x"dd",x"87"),
   860 => (x"c4",x"86",x"70",x"98"),
   861 => (x"05",x"c5",x"87",x"c0"),
   862 => (x"48",x"c1",x"c0",x"87"),
   863 => (x"c1",x"84",x"c1",x"cc"),
   864 => (x"ee",x"bf",x"49",x"74"),
   865 => (x"99",x"05",x"cc",x"87"),
   866 => (x"c1",x"cd",x"ee",x"bf"),
   867 => (x"49",x"f6",x"f1",x"87"),
   868 => (x"c1",x"cd",x"f2",x"58"),
   869 => (x"d4",x"66",x"48",x"c8"),
   870 => (x"c0",x"80",x"d8",x"a6"),
   871 => (x"58",x"c1",x"85",x"6e"),
   872 => (x"b7",x"ad",x"04",x"fe"),
   873 => (x"e4",x"87",x"cf",x"87"),
   874 => (x"73",x"1e",x"c0",x"ec"),
   875 => (x"f2",x"1e",x"cb",x"f6"),
   876 => (x"87",x"c8",x"86",x"c0"),
   877 => (x"48",x"c5",x"87",x"c1"),
   878 => (x"cd",x"ea",x"bf",x"48"),
   879 => (x"26",x"e5",x"da",x"87"),
   880 => (x"1e",x"f3",x"09",x"97"),
   881 => (x"79",x"09",x"71",x"48"),
   882 => (x"26",x"4f",x"0e",x"5e"),
   883 => (x"5b",x"5c",x"0e",x"71"),
   884 => (x"4b",x"c0",x"4c",x"13"),
   885 => (x"4a",x"72",x"9a",x"02"),
   886 => (x"cd",x"87",x"72",x"49"),
   887 => (x"e2",x"87",x"c1",x"84"),
   888 => (x"13",x"4a",x"72",x"9a"),
   889 => (x"05",x"f3",x"87",x"74"),
   890 => (x"48",x"c2",x"87",x"26"),
   891 => (x"4d",x"26",x"4c",x"26"),
   892 => (x"4b",x"26",x"4f",x"0e"),
   893 => (x"5e",x"5b",x"5c",x"5d"),
   894 => (x"0e",x"fc",x"86",x"71"),
   895 => (x"4a",x"c0",x"e0",x"66"),
   896 => (x"4c",x"c1",x"cd",x"f2"),
   897 => (x"4b",x"c0",x"7e",x"72"),
   898 => (x"9a",x"05",x"ce",x"87"),
   899 => (x"c1",x"cd",x"f3",x"4b"),
   900 => (x"c1",x"cd",x"f2",x"48"),
   901 => (x"c0",x"f0",x"50",x"c1"),
   902 => (x"d2",x"87",x"72",x"9a"),
   903 => (x"02",x"c0",x"e9",x"87"),
   904 => (x"d4",x"66",x"4d",x"72"),
   905 => (x"1e",x"72",x"49",x"75"),
   906 => (x"4a",x"ca",x"cf",x"87"),
   907 => (x"26",x"4a",x"c0",x"fa"),
   908 => (x"dd",x"81",x"11",x"53"),
   909 => (x"71",x"1e",x"72",x"49"),
   910 => (x"75",x"4a",x"c9",x"fe"),
   911 => (x"87",x"70",x"4a",x"26"),
   912 => (x"49",x"c1",x"8c",x"72"),
   913 => (x"9a",x"05",x"ff",x"da"),
   914 => (x"87",x"c0",x"b7",x"ac"),
   915 => (x"06",x"dd",x"87",x"c0"),
   916 => (x"e4",x"66",x"02",x"c5"),
   917 => (x"87",x"c0",x"f0",x"4a"),
   918 => (x"c3",x"87",x"c0",x"e0"),
   919 => (x"4a",x"73",x"0a",x"97"),
   920 => (x"7a",x"0a",x"c1",x"83"),
   921 => (x"8c",x"c0",x"b7",x"ac"),
   922 => (x"01",x"ff",x"e3",x"87"),
   923 => (x"c1",x"cd",x"f2",x"ab"),
   924 => (x"02",x"de",x"87",x"d8"),
   925 => (x"66",x"4c",x"dc",x"66"),
   926 => (x"1e",x"c1",x"8b",x"97"),
   927 => (x"6b",x"49",x"74",x"0f"),
   928 => (x"c4",x"86",x"6e",x"48"),
   929 => (x"c1",x"80",x"c4",x"a6"),
   930 => (x"58",x"c1",x"cd",x"f2"),
   931 => (x"ab",x"05",x"ff",x"e5"),
   932 => (x"87",x"6e",x"48",x"fc"),
   933 => (x"8e",x"26",x"4d",x"26"),
   934 => (x"4c",x"26",x"4b",x"26"),
   935 => (x"4f",x"30",x"31",x"32"),
   936 => (x"33",x"34",x"35",x"36"),
   937 => (x"37",x"38",x"39",x"41"),
   938 => (x"42",x"43",x"44",x"45"),
   939 => (x"46",x"00",x"0e",x"5e"),
   940 => (x"5b",x"5c",x"5d",x"0e"),
   941 => (x"71",x"4b",x"ff",x"4d"),
   942 => (x"13",x"4c",x"74",x"9c"),
   943 => (x"02",x"d8",x"87",x"c1"),
   944 => (x"85",x"d4",x"66",x"1e"),
   945 => (x"74",x"49",x"d4",x"66"),
   946 => (x"0f",x"c4",x"86",x"74"),
   947 => (x"a8",x"05",x"c7",x"87"),
   948 => (x"13",x"4c",x"74",x"9c"),
   949 => (x"05",x"e8",x"87",x"75"),
   950 => (x"48",x"26",x"4d",x"26"),
   951 => (x"4c",x"26",x"4b",x"26"),
   952 => (x"4f",x"0e",x"5e",x"5b"),
   953 => (x"5c",x"5d",x"0e",x"e8"),
   954 => (x"86",x"c4",x"a6",x"59"),
   955 => (x"c0",x"e8",x"66",x"4d"),
   956 => (x"c0",x"4c",x"c8",x"a6"),
   957 => (x"48",x"c0",x"78",x"6e"),
   958 => (x"97",x"bf",x"4b",x"6e"),
   959 => (x"48",x"c1",x"80",x"c4"),
   960 => (x"a6",x"58",x"73",x"9b"),
   961 => (x"02",x"c6",x"d3",x"87"),
   962 => (x"c8",x"66",x"02",x"c5"),
   963 => (x"db",x"87",x"cc",x"a6"),
   964 => (x"48",x"c0",x"78",x"fc"),
   965 => (x"80",x"c0",x"78",x"73"),
   966 => (x"4a",x"c0",x"e0",x"8a"),
   967 => (x"02",x"c3",x"c6",x"87"),
   968 => (x"c3",x"8a",x"02",x"c3"),
   969 => (x"c0",x"87",x"c2",x"8a"),
   970 => (x"02",x"c2",x"e8",x"87"),
   971 => (x"c2",x"8a",x"02",x"c2"),
   972 => (x"f4",x"87",x"c4",x"8a"),
   973 => (x"02",x"c2",x"ee",x"87"),
   974 => (x"c2",x"8a",x"02",x"c2"),
   975 => (x"e8",x"87",x"c3",x"8a"),
   976 => (x"02",x"c2",x"ea",x"87"),
   977 => (x"d4",x"8a",x"02",x"c0"),
   978 => (x"f6",x"87",x"d4",x"8a"),
   979 => (x"02",x"c1",x"c0",x"87"),
   980 => (x"ca",x"8a",x"02",x"c0"),
   981 => (x"f2",x"87",x"c1",x"8a"),
   982 => (x"02",x"c1",x"e1",x"87"),
   983 => (x"c1",x"8a",x"02",x"df"),
   984 => (x"87",x"c8",x"8a",x"02"),
   985 => (x"c1",x"ce",x"87",x"c4"),
   986 => (x"8a",x"02",x"c0",x"e3"),
   987 => (x"87",x"c3",x"8a",x"02"),
   988 => (x"c0",x"e5",x"87",x"c2"),
   989 => (x"8a",x"02",x"c8",x"87"),
   990 => (x"c3",x"8a",x"02",x"d3"),
   991 => (x"87",x"c1",x"fa",x"87"),
   992 => (x"cc",x"a6",x"48",x"ca"),
   993 => (x"78",x"c2",x"d2",x"87"),
   994 => (x"cc",x"a6",x"48",x"c2"),
   995 => (x"78",x"c2",x"ca",x"87"),
   996 => (x"cc",x"a6",x"48",x"d0"),
   997 => (x"78",x"c2",x"c2",x"87"),
   998 => (x"c0",x"f0",x"66",x"1e"),
   999 => (x"c0",x"f0",x"66",x"1e"),
  1000 => (x"c4",x"85",x"75",x"4a"),
  1001 => (x"c4",x"8a",x"6a",x"49"),
  1002 => (x"fc",x"c3",x"87",x"c8"),
  1003 => (x"86",x"70",x"49",x"71"),
  1004 => (x"a4",x"4c",x"c1",x"e5"),
  1005 => (x"87",x"c8",x"a6",x"48"),
  1006 => (x"c1",x"78",x"c1",x"dd"),
  1007 => (x"87",x"c0",x"f0",x"66"),
  1008 => (x"1e",x"c4",x"85",x"75"),
  1009 => (x"4a",x"c4",x"8a",x"6a"),
  1010 => (x"49",x"c0",x"f0",x"66"),
  1011 => (x"0f",x"c4",x"86",x"c1"),
  1012 => (x"84",x"c1",x"c6",x"87"),
  1013 => (x"c0",x"f0",x"66",x"1e"),
  1014 => (x"c0",x"e5",x"49",x"c0"),
  1015 => (x"f0",x"66",x"0f",x"c4"),
  1016 => (x"86",x"c1",x"84",x"c0"),
  1017 => (x"f4",x"87",x"c8",x"a6"),
  1018 => (x"48",x"c1",x"78",x"c0"),
  1019 => (x"ec",x"87",x"d0",x"a6"),
  1020 => (x"48",x"c1",x"78",x"f8"),
  1021 => (x"80",x"c1",x"78",x"c0"),
  1022 => (x"e0",x"87",x"c0",x"f0"),
  1023 => (x"ab",x"06",x"da",x"87"),
  1024 => (x"c0",x"f9",x"ab",x"03"),
  1025 => (x"d4",x"87",x"d4",x"66"),
  1026 => (x"49",x"ca",x"91",x"73"),
  1027 => (x"4a",x"c0",x"f0",x"8a"),
  1028 => (x"d4",x"a6",x"48",x"72"),
  1029 => (x"a1",x"78",x"f4",x"80"),
  1030 => (x"c1",x"78",x"cc",x"66"),
  1031 => (x"02",x"c1",x"ea",x"87"),
  1032 => (x"c4",x"85",x"75",x"49"),
  1033 => (x"c4",x"89",x"a6",x"48"),
  1034 => (x"69",x"78",x"c1",x"e4"),
  1035 => (x"ab",x"05",x"d8",x"87"),
  1036 => (x"c4",x"66",x"48",x"c0"),
  1037 => (x"b7",x"a8",x"03",x"cf"),
  1038 => (x"87",x"c0",x"ed",x"49"),
  1039 => (x"f6",x"c1",x"87",x"c4"),
  1040 => (x"66",x"48",x"c0",x"08"),
  1041 => (x"88",x"c8",x"a6",x"58"),
  1042 => (x"d0",x"66",x"1e",x"d8"),
  1043 => (x"66",x"1e",x"c0",x"f8"),
  1044 => (x"66",x"1e",x"c0",x"f8"),
  1045 => (x"66",x"1e",x"dc",x"66"),
  1046 => (x"1e",x"d8",x"66",x"49"),
  1047 => (x"f6",x"d4",x"87",x"d4"),
  1048 => (x"86",x"70",x"49",x"71"),
  1049 => (x"a4",x"4c",x"c0",x"e1"),
  1050 => (x"87",x"c0",x"e5",x"ab"),
  1051 => (x"05",x"cf",x"87",x"d0"),
  1052 => (x"a6",x"48",x"c0",x"78"),
  1053 => (x"c4",x"80",x"c0",x"78"),
  1054 => (x"f4",x"80",x"c1",x"78"),
  1055 => (x"cc",x"87",x"c0",x"f0"),
  1056 => (x"66",x"1e",x"73",x"49"),
  1057 => (x"c0",x"f0",x"66",x"0f"),
  1058 => (x"c4",x"86",x"6e",x"97"),
  1059 => (x"bf",x"4b",x"6e",x"48"),
  1060 => (x"c1",x"80",x"c4",x"a6"),
  1061 => (x"58",x"73",x"9b",x"05"),
  1062 => (x"f9",x"ed",x"87",x"74"),
  1063 => (x"48",x"e8",x"8e",x"26"),
  1064 => (x"4d",x"26",x"4c",x"26"),
  1065 => (x"4b",x"26",x"4f",x"1e"),
  1066 => (x"c0",x"1e",x"c0",x"f7"),
  1067 => (x"c0",x"1e",x"d0",x"a6"),
  1068 => (x"1e",x"d0",x"66",x"49"),
  1069 => (x"f8",x"ea",x"87",x"f4"),
  1070 => (x"8e",x"26",x"4f",x"1e"),
  1071 => (x"73",x"1e",x"72",x"9a"),
  1072 => (x"02",x"c0",x"e7",x"87"),
  1073 => (x"c0",x"48",x"c1",x"4b"),
  1074 => (x"72",x"a9",x"06",x"d1"),
  1075 => (x"87",x"72",x"82",x"06"),
  1076 => (x"c9",x"87",x"73",x"83"),
  1077 => (x"72",x"a9",x"01",x"f4"),
  1078 => (x"87",x"c3",x"87",x"c1"),
  1079 => (x"b2",x"3a",x"72",x"a9"),
  1080 => (x"03",x"89",x"73",x"80"),
  1081 => (x"07",x"c1",x"2a",x"2b"),
  1082 => (x"05",x"f3",x"87",x"26"),
  1083 => (x"4b",x"26",x"4f",x"1e"),
  1084 => (x"75",x"1e",x"c4",x"4d"),
  1085 => (x"71",x"b7",x"a1",x"04"),
  1086 => (x"ff",x"b9",x"c1",x"81"),
  1087 => (x"c3",x"bd",x"07",x"72"),
  1088 => (x"b7",x"a2",x"04",x"ff"),
  1089 => (x"ba",x"c1",x"82",x"c1"),
  1090 => (x"bd",x"07",x"fe",x"ee"),
  1091 => (x"87",x"c1",x"2d",x"04"),
  1092 => (x"ff",x"b8",x"c1",x"80"),
  1093 => (x"07",x"2d",x"04",x"ff"),
  1094 => (x"b9",x"c1",x"81",x"07"),
  1095 => (x"26",x"4d",x"26",x"4f"),
	others => (others => x"00")
);

-- Xilinx XST attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "no_rw_check";

-- Altera Quartus attributes
attribute ramstyle: string;
attribute ramstyle of ram: signal is "no_rw_check";

signal q_local : word_t;

begin
    
	process(clk,q_local)
	begin

		q(31 downto 24)<=q_local(0);
		q(23 downto 16)<=q_local(1);
		q(15 downto 8)<=q_local(2);
		q(7 downto 0)<=q_local(3);

		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel(3) = '1') then
					ram(to_integer(unsigned(addr)))(3) <= d(7 downto 0);
				end if;
				if bytesel(2) = '1' then
					ram(to_integer(unsigned(addr)))(2) <= d(15 downto 8);
				end if;
				if bytesel(1) = '1' then
					ram(to_integer(unsigned(addr)))(1) <= d(23 downto 16);
				end if;
				if bytesel(0) = '1' then
					ram(to_integer(unsigned(addr)))(0) <= d(31 downto 24);
				end if;
			end if;
			q_local <= ram(to_integer(unsigned(addr)));
		end if;
	end process;

end arch;

