library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM-2 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
type ram_type is array (0 to 2 ** (maxAddrBitBRAM-3) - 1) of word_t;

signal ram : ram_type :=
(
     0 => (x"01",x"da",x"87",x"04"),
     1 => (x"dd",x"87",x"0e",x"58"),
     2 => (x"5e",x"59",x"5a",x"0e"),
     3 => (x"27",x"00",x"00",x"00"),
     4 => (x"2c",x"0f",x"26",x"4a"),
     5 => (x"26",x"49",x"26",x"48"),
     6 => (x"ff",x"80",x"26",x"08"),
     7 => (x"4f",x"27",x"00",x"00"),
     8 => (x"00",x"2d",x"4f",x"27"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"4f",x"00",x"fd",x"87"),
    11 => (x"4f",x"c1",x"ce",x"e4"),
    12 => (x"4e",x"c9",x"c0",x"86"),
    13 => (x"c1",x"ce",x"e4",x"49"),
    14 => (x"c1",x"c5",x"c0",x"48"),
    15 => (x"89",x"d0",x"89",x"03"),
    16 => (x"c0",x"40",x"40",x"40"),
    17 => (x"40",x"f6",x"87",x"d0"),
    18 => (x"81",x"05",x"c0",x"50"),
    19 => (x"c1",x"89",x"05",x"f9"),
    20 => (x"87",x"c1",x"c4",x"fd"),
    21 => (x"4d",x"c1",x"c4",x"fd"),
    22 => (x"4c",x"74",x"ad",x"02"),
    23 => (x"c4",x"87",x"24",x"0f"),
    24 => (x"f7",x"87",x"c2",x"da"),
    25 => (x"87",x"c1",x"c4",x"fd"),
    26 => (x"4d",x"c1",x"c4",x"fd"),
    27 => (x"4c",x"74",x"ad",x"02"),
    28 => (x"c6",x"87",x"c4",x"8c"),
    29 => (x"6c",x"0f",x"f5",x"87"),
    30 => (x"00",x"fd",x"87",x"0e"),
    31 => (x"5e",x"5b",x"5c",x"0e"),
    32 => (x"c0",x"e8",x"c0",x"c0"),
    33 => (x"c0",x"4b",x"c9",x"e2"),
    34 => (x"4c",x"c9",x"f4",x"bf"),
    35 => (x"4a",x"c1",x"8a",x"02"),
    36 => (x"cb",x"87",x"74",x"49"),
    37 => (x"c1",x"84",x"11",x"53"),
    38 => (x"c1",x"8a",x"05",x"f5"),
    39 => (x"87",x"c2",x"87",x"26"),
    40 => (x"4d",x"26",x"4c",x"26"),
    41 => (x"4b",x"26",x"4f",x"0e"),
    42 => (x"5e",x"5b",x"5c",x"0e"),
    43 => (x"71",x"4b",x"c0",x"e8"),
    44 => (x"c0",x"c0",x"c0",x"4c"),
    45 => (x"e7",x"48",x"c0",x"e0"),
    46 => (x"50",x"e3",x"48",x"c8"),
    47 => (x"50",x"e3",x"48",x"c6"),
    48 => (x"50",x"e7",x"48",x"c0"),
    49 => (x"e1",x"50",x"73",x"4a"),
    50 => (x"c8",x"b7",x"2a",x"ca"),
    51 => (x"a4",x"49",x"71",x"0a"),
    52 => (x"97",x"7a",x"73",x"4a"),
    53 => (x"c3",x"ff",x"9a",x"cb"),
    54 => (x"a4",x"49",x"71",x"0a"),
    55 => (x"97",x"7a",x"e7",x"48"),
    56 => (x"c0",x"e0",x"50",x"e3"),
    57 => (x"48",x"c8",x"50",x"e3"),
    58 => (x"48",x"c0",x"50",x"e7"),
    59 => (x"48",x"c0",x"e1",x"50"),
    60 => (x"fe",x"ee",x"87",x"1e"),
    61 => (x"73",x"1e",x"c2",x"c0"),
    62 => (x"c0",x"4b",x"73",x"0f"),
    63 => (x"fe",x"e4",x"87",x"1e"),
    64 => (x"73",x"1e",x"eb",x"48"),
    65 => (x"c3",x"ef",x"50",x"e7"),
    66 => (x"48",x"c0",x"e0",x"50"),
    67 => (x"e3",x"48",x"c8",x"50"),
    68 => (x"e3",x"48",x"c6",x"50"),
    69 => (x"e7",x"48",x"c0",x"e1"),
    70 => (x"50",x"ff",x"c2",x"48"),
    71 => (x"c1",x"9f",x"78",x"e7"),
    72 => (x"48",x"c0",x"e0",x"50"),
    73 => (x"e3",x"48",x"c4",x"50"),
    74 => (x"e3",x"48",x"c2",x"50"),
    75 => (x"e7",x"48",x"c0",x"e1"),
    76 => (x"50",x"e7",x"48",x"c0"),
    77 => (x"e0",x"50",x"e3",x"48"),
    78 => (x"c8",x"50",x"e3",x"48"),
    79 => (x"c7",x"50",x"e7",x"48"),
    80 => (x"c0",x"e1",x"50",x"fc"),
    81 => (x"f5",x"87",x"c0",x"ff"),
    82 => (x"ff",x"49",x"fd",x"da"),
    83 => (x"87",x"c0",x"fc",x"c0"),
    84 => (x"4b",x"c8",x"ee",x"49"),
    85 => (x"c0",x"f2",x"cf",x"87"),
    86 => (x"d1",x"dd",x"87",x"70"),
    87 => (x"98",x"02",x"c1",x"cb"),
    88 => (x"87",x"c0",x"ff",x"f0"),
    89 => (x"4b",x"c8",x"d7",x"49"),
    90 => (x"c0",x"f1",x"fb",x"87"),
    91 => (x"d7",x"d0",x"87",x"70"),
    92 => (x"98",x"02",x"c0",x"e7"),
    93 => (x"87",x"c3",x"f0",x"4b"),
    94 => (x"c2",x"c0",x"c0",x"1e"),
    95 => (x"c6",x"fe",x"49",x"c0"),
    96 => (x"ee",x"f1",x"87",x"c4"),
    97 => (x"86",x"70",x"98",x"02"),
    98 => (x"c9",x"87",x"c3",x"ff"),
    99 => (x"4b",x"fd",x"e3",x"87"),
   100 => (x"c0",x"e0",x"87",x"c7"),
   101 => (x"ca",x"49",x"c0",x"f1"),
   102 => (x"cd",x"87",x"d7",x"87"),
   103 => (x"c7",x"df",x"49",x"c0"),
   104 => (x"f1",x"c4",x"87",x"c7"),
   105 => (x"fb",x"49",x"c0",x"f0"),
   106 => (x"fd",x"87",x"c7",x"87"),
   107 => (x"c9",x"c4",x"49",x"c0"),
   108 => (x"f0",x"f4",x"87",x"73"),
   109 => (x"49",x"fb",x"ef",x"87"),
   110 => (x"fe",x"d2",x"87",x"fb"),
   111 => (x"e5",x"87",x"38",x"33"),
   112 => (x"32",x"4f",x"53",x"44"),
   113 => (x"41",x"42",x"42",x"49"),
   114 => (x"4e",x"00",x"43",x"61"),
   115 => (x"6e",x"27",x"74",x"20"),
   116 => (x"6c",x"6f",x"61",x"64"),
   117 => (x"20",x"66",x"69",x"72"),
   118 => (x"6d",x"77",x"61",x"72"),
   119 => (x"65",x"0a",x"00",x"55"),
   120 => (x"6e",x"61",x"62",x"6c"),
   121 => (x"65",x"20",x"74",x"6f"),
   122 => (x"20",x"6c",x"6f",x"63"),
   123 => (x"61",x"74",x"65",x"20"),
   124 => (x"70",x"61",x"72",x"74"),
   125 => (x"69",x"74",x"69",x"6f"),
   126 => (x"6e",x"0a",x"00",x"55"),
   127 => (x"6e",x"61",x"62",x"6c"),
   128 => (x"65",x"20",x"74",x"6f"),
   129 => (x"20",x"6c",x"6f",x"63"),
   130 => (x"61",x"74",x"65",x"20"),
   131 => (x"70",x"61",x"72",x"74"),
   132 => (x"69",x"74",x"69",x"6f"),
   133 => (x"6e",x"0a",x"00",x"48"),
   134 => (x"75",x"6e",x"74",x"69"),
   135 => (x"6e",x"67",x"20",x"66"),
   136 => (x"6f",x"72",x"20",x"70"),
   137 => (x"61",x"72",x"74",x"69"),
   138 => (x"74",x"69",x"6f",x"6e"),
   139 => (x"0a",x"00",x"49",x"6e"),
   140 => (x"69",x"74",x"69",x"61"),
   141 => (x"6c",x"69",x"7a",x"69"),
   142 => (x"6e",x"67",x"20",x"53"),
   143 => (x"44",x"20",x"63",x"61"),
   144 => (x"72",x"64",x"0a",x"00"),
   145 => (x"46",x"61",x"69",x"6c"),
   146 => (x"65",x"64",x"20",x"74"),
   147 => (x"6f",x"20",x"69",x"6e"),
   148 => (x"69",x"74",x"69",x"61"),
   149 => (x"6c",x"69",x"7a",x"65"),
   150 => (x"20",x"53",x"44",x"20"),
   151 => (x"63",x"61",x"72",x"64"),
   152 => (x"0a",x"00",x"00",x"00"),
   153 => (x"00",x"00",x"00",x"00"),
   154 => (x"00",x"08",x"33",x"fc"),
   155 => (x"0f",x"ff",x"00",x"df"),
   156 => (x"f1",x"80",x"60",x"f6"),
   157 => (x"00",x"00",x"00",x"12"),
   158 => (x"1e",x"e4",x"86",x"e3"),
   159 => (x"48",x"c3",x"ff",x"50"),
   160 => (x"e3",x"97",x"bf",x"48"),
   161 => (x"c4",x"a6",x"58",x"6e"),
   162 => (x"49",x"c3",x"ff",x"99"),
   163 => (x"e3",x"48",x"c3",x"ff"),
   164 => (x"50",x"c8",x"31",x"e3"),
   165 => (x"97",x"bf",x"48",x"c8"),
   166 => (x"a6",x"58",x"c4",x"66"),
   167 => (x"48",x"c3",x"ff",x"98"),
   168 => (x"cc",x"a6",x"58",x"c8"),
   169 => (x"66",x"b1",x"e3",x"48"),
   170 => (x"c3",x"ff",x"50",x"c8"),
   171 => (x"31",x"e3",x"97",x"bf"),
   172 => (x"48",x"d0",x"a6",x"58"),
   173 => (x"cc",x"66",x"48",x"c3"),
   174 => (x"ff",x"98",x"d4",x"a6"),
   175 => (x"58",x"d0",x"66",x"b1"),
   176 => (x"e3",x"48",x"c3",x"ff"),
   177 => (x"50",x"c8",x"31",x"e3"),
   178 => (x"97",x"bf",x"48",x"d8"),
   179 => (x"a6",x"58",x"d4",x"66"),
   180 => (x"48",x"c3",x"ff",x"98"),
   181 => (x"dc",x"a6",x"58",x"d8"),
   182 => (x"66",x"b1",x"71",x"48"),
   183 => (x"e4",x"8e",x"26",x"4f"),
   184 => (x"0e",x"5e",x"5b",x"5c"),
   185 => (x"0e",x"1e",x"71",x"4a"),
   186 => (x"72",x"49",x"c3",x"ff"),
   187 => (x"99",x"e3",x"09",x"97"),
   188 => (x"79",x"09",x"c1",x"c5"),
   189 => (x"c0",x"bf",x"05",x"c8"),
   190 => (x"87",x"d0",x"66",x"48"),
   191 => (x"c9",x"30",x"d4",x"a6"),
   192 => (x"58",x"d0",x"66",x"49"),
   193 => (x"d8",x"29",x"c3",x"ff"),
   194 => (x"99",x"e3",x"09",x"97"),
   195 => (x"79",x"09",x"d0",x"66"),
   196 => (x"49",x"d0",x"29",x"c3"),
   197 => (x"ff",x"99",x"e3",x"09"),
   198 => (x"97",x"79",x"09",x"d0"),
   199 => (x"66",x"49",x"c8",x"29"),
   200 => (x"c3",x"ff",x"99",x"e3"),
   201 => (x"09",x"97",x"79",x"09"),
   202 => (x"d0",x"66",x"49",x"c3"),
   203 => (x"ff",x"99",x"e3",x"09"),
   204 => (x"97",x"79",x"09",x"72"),
   205 => (x"49",x"d0",x"29",x"c3"),
   206 => (x"ff",x"99",x"e3",x"09"),
   207 => (x"97",x"79",x"09",x"97"),
   208 => (x"bf",x"48",x"c4",x"a6"),
   209 => (x"58",x"6e",x"4b",x"c3"),
   210 => (x"ff",x"9b",x"c9",x"f0"),
   211 => (x"ff",x"4c",x"c3",x"ff"),
   212 => (x"ab",x"05",x"dc",x"87"),
   213 => (x"e3",x"48",x"c3",x"ff"),
   214 => (x"50",x"e3",x"97",x"bf"),
   215 => (x"48",x"c4",x"a6",x"58"),
   216 => (x"6e",x"4b",x"c3",x"ff"),
   217 => (x"9b",x"c1",x"8c",x"02"),
   218 => (x"c6",x"87",x"c3",x"ff"),
   219 => (x"ab",x"02",x"e4",x"87"),
   220 => (x"73",x"4a",x"c4",x"b7"),
   221 => (x"2a",x"c0",x"f0",x"a2"),
   222 => (x"49",x"c0",x"e9",x"e0"),
   223 => (x"87",x"73",x"4a",x"cf"),
   224 => (x"9a",x"c0",x"f0",x"a2"),
   225 => (x"49",x"c0",x"e9",x"d4"),
   226 => (x"87",x"73",x"48",x"26"),
   227 => (x"c2",x"87",x"26",x"4d"),
   228 => (x"26",x"4c",x"26",x"4b"),
   229 => (x"26",x"4f",x"1e",x"c0"),
   230 => (x"49",x"e3",x"48",x"c3"),
   231 => (x"ff",x"50",x"c1",x"81"),
   232 => (x"c3",x"c8",x"b7",x"a9"),
   233 => (x"04",x"f2",x"87",x"26"),
   234 => (x"4f",x"1e",x"73",x"1e"),
   235 => (x"e8",x"87",x"c4",x"f8"),
   236 => (x"df",x"4b",x"c0",x"1e"),
   237 => (x"c0",x"ff",x"f0",x"c1"),
   238 => (x"f7",x"49",x"fc",x"e3"),
   239 => (x"87",x"c4",x"86",x"c1"),
   240 => (x"a8",x"05",x"c0",x"e8"),
   241 => (x"87",x"e3",x"48",x"c3"),
   242 => (x"ff",x"50",x"c1",x"c0"),
   243 => (x"c0",x"c0",x"c0",x"c0"),
   244 => (x"1e",x"c0",x"e1",x"f0"),
   245 => (x"c1",x"e9",x"49",x"fc"),
   246 => (x"c6",x"87",x"c4",x"86"),
   247 => (x"70",x"98",x"05",x"c9"),
   248 => (x"87",x"e3",x"48",x"c3"),
   249 => (x"ff",x"50",x"c1",x"48"),
   250 => (x"cb",x"87",x"fe",x"e9"),
   251 => (x"87",x"c1",x"8b",x"05"),
   252 => (x"fe",x"ff",x"87",x"c0"),
   253 => (x"48",x"fe",x"da",x"87"),
   254 => (x"43",x"4d",x"44",x"34"),
   255 => (x"31",x"20",x"25",x"64"),
   256 => (x"0a",x"00",x"43",x"4d"),
   257 => (x"44",x"35",x"35",x"20"),
   258 => (x"25",x"64",x"0a",x"00"),
   259 => (x"43",x"4d",x"44",x"34"),
   260 => (x"31",x"20",x"25",x"64"),
   261 => (x"0a",x"00",x"43",x"4d"),
   262 => (x"44",x"35",x"35",x"20"),
   263 => (x"25",x"64",x"0a",x"00"),
   264 => (x"69",x"6e",x"69",x"74"),
   265 => (x"20",x"25",x"64",x"0a"),
   266 => (x"20",x"20",x"00",x"69"),
   267 => (x"6e",x"69",x"74",x"20"),
   268 => (x"25",x"64",x"0a",x"20"),
   269 => (x"20",x"00",x"43",x"6d"),
   270 => (x"64",x"5f",x"69",x"6e"),
   271 => (x"69",x"74",x"0a",x"00"),
   272 => (x"43",x"4d",x"44",x"38"),
   273 => (x"5f",x"34",x"20",x"72"),
   274 => (x"65",x"73",x"70",x"6f"),
   275 => (x"6e",x"73",x"65",x"3a"),
   276 => (x"20",x"25",x"64",x"0a"),
   277 => (x"00",x"43",x"4d",x"44"),
   278 => (x"35",x"38",x"20",x"25"),
   279 => (x"64",x"0a",x"20",x"20"),
   280 => (x"00",x"43",x"4d",x"44"),
   281 => (x"35",x"38",x"5f",x"32"),
   282 => (x"20",x"25",x"64",x"0a"),
   283 => (x"20",x"20",x"00",x"43"),
   284 => (x"4d",x"44",x"35",x"38"),
   285 => (x"20",x"25",x"64",x"0a"),
   286 => (x"20",x"20",x"00",x"53"),
   287 => (x"44",x"48",x"43",x"20"),
   288 => (x"49",x"6e",x"69",x"74"),
   289 => (x"69",x"61",x"6c",x"69"),
   290 => (x"7a",x"61",x"74",x"69"),
   291 => (x"6f",x"6e",x"20",x"65"),
   292 => (x"72",x"72",x"6f",x"72"),
   293 => (x"21",x"0a",x"00",x"63"),
   294 => (x"6d",x"64",x"5f",x"43"),
   295 => (x"4d",x"44",x"38",x"20"),
   296 => (x"72",x"65",x"73",x"70"),
   297 => (x"6f",x"6e",x"73",x"65"),
   298 => (x"3a",x"20",x"25",x"64"),
   299 => (x"0a",x"00",x"52",x"65"),
   300 => (x"61",x"64",x"20",x"63"),
   301 => (x"6f",x"6d",x"6d",x"61"),
   302 => (x"6e",x"64",x"20",x"66"),
   303 => (x"61",x"69",x"6c",x"65"),
   304 => (x"64",x"20",x"61",x"74"),
   305 => (x"20",x"25",x"64",x"20"),
   306 => (x"28",x"25",x"64",x"29"),
   307 => (x"0a",x"00",x"1e",x"73"),
   308 => (x"1e",x"e3",x"48",x"c3"),
   309 => (x"ff",x"50",x"d0",x"f6"),
   310 => (x"49",x"c0",x"e4",x"ca"),
   311 => (x"87",x"d3",x"4b",x"c0"),
   312 => (x"1e",x"c0",x"ff",x"f0"),
   313 => (x"c1",x"c1",x"49",x"f7"),
   314 => (x"f6",x"87",x"c4",x"86"),
   315 => (x"70",x"98",x"05",x"c9"),
   316 => (x"87",x"e3",x"48",x"c3"),
   317 => (x"ff",x"50",x"c1",x"48"),
   318 => (x"cb",x"87",x"fa",x"d9"),
   319 => (x"87",x"c1",x"8b",x"05"),
   320 => (x"ff",x"dc",x"87",x"c0"),
   321 => (x"48",x"fa",x"ca",x"87"),
   322 => (x"1e",x"73",x"1e",x"1e"),
   323 => (x"fa",x"c7",x"87",x"c6"),
   324 => (x"ea",x"1e",x"c0",x"e1"),
   325 => (x"f0",x"c1",x"c8",x"49"),
   326 => (x"f7",x"c5",x"87",x"70"),
   327 => (x"4b",x"73",x"1e",x"d2"),
   328 => (x"d7",x"49",x"c0",x"ee"),
   329 => (x"de",x"87",x"c8",x"86"),
   330 => (x"c1",x"ab",x"02",x"c8"),
   331 => (x"87",x"fe",x"de",x"87"),
   332 => (x"c0",x"48",x"c1",x"ff"),
   333 => (x"87",x"f5",x"c0",x"87"),
   334 => (x"70",x"49",x"cf",x"ff"),
   335 => (x"ff",x"99",x"c6",x"ea"),
   336 => (x"a9",x"02",x"c8",x"87"),
   337 => (x"fe",x"c7",x"87",x"c0"),
   338 => (x"48",x"c1",x"e8",x"87"),
   339 => (x"e3",x"48",x"c3",x"ff"),
   340 => (x"50",x"c0",x"f1",x"4b"),
   341 => (x"f9",x"d2",x"87",x"70"),
   342 => (x"98",x"02",x"c1",x"c6"),
   343 => (x"87",x"c0",x"1e",x"c0"),
   344 => (x"ff",x"f0",x"c1",x"fa"),
   345 => (x"49",x"f5",x"f8",x"87"),
   346 => (x"c4",x"86",x"70",x"98"),
   347 => (x"05",x"c0",x"f3",x"87"),
   348 => (x"e3",x"48",x"c3",x"ff"),
   349 => (x"50",x"e3",x"97",x"bf"),
   350 => (x"48",x"c4",x"a6",x"58"),
   351 => (x"6e",x"49",x"c3",x"ff"),
   352 => (x"99",x"e3",x"48",x"c3"),
   353 => (x"ff",x"50",x"e3",x"48"),
   354 => (x"c3",x"ff",x"50",x"e3"),
   355 => (x"48",x"c3",x"ff",x"50"),
   356 => (x"e3",x"48",x"c3",x"ff"),
   357 => (x"50",x"c1",x"c0",x"99"),
   358 => (x"02",x"c4",x"87",x"c1"),
   359 => (x"48",x"d5",x"87",x"c0"),
   360 => (x"48",x"d1",x"87",x"c2"),
   361 => (x"ab",x"05",x"c4",x"87"),
   362 => (x"c0",x"48",x"c8",x"87"),
   363 => (x"c1",x"8b",x"05",x"fe"),
   364 => (x"e2",x"87",x"c0",x"48"),
   365 => (x"26",x"f7",x"da",x"87"),
   366 => (x"1e",x"73",x"1e",x"c1"),
   367 => (x"c5",x"c0",x"48",x"c1"),
   368 => (x"78",x"eb",x"48",x"c3"),
   369 => (x"ef",x"50",x"c7",x"4b"),
   370 => (x"e7",x"48",x"c3",x"50"),
   371 => (x"f7",x"c7",x"87",x"e7"),
   372 => (x"48",x"c2",x"50",x"e3"),
   373 => (x"48",x"c3",x"ff",x"50"),
   374 => (x"c0",x"1e",x"c0",x"e5"),
   375 => (x"d0",x"c1",x"c0",x"49"),
   376 => (x"f3",x"fd",x"87",x"c4"),
   377 => (x"86",x"c1",x"a8",x"05"),
   378 => (x"c2",x"87",x"c1",x"4b"),
   379 => (x"c2",x"ab",x"05",x"c5"),
   380 => (x"87",x"c0",x"48",x"c0"),
   381 => (x"f1",x"87",x"c1",x"8b"),
   382 => (x"05",x"ff",x"cc",x"87"),
   383 => (x"fc",x"c9",x"87",x"c1"),
   384 => (x"c5",x"c4",x"58",x"c1"),
   385 => (x"c5",x"c0",x"bf",x"05"),
   386 => (x"cd",x"87",x"c1",x"1e"),
   387 => (x"c0",x"ff",x"f0",x"c1"),
   388 => (x"d0",x"49",x"f3",x"cb"),
   389 => (x"87",x"c4",x"86",x"e3"),
   390 => (x"48",x"c3",x"ff",x"50"),
   391 => (x"e7",x"48",x"c3",x"50"),
   392 => (x"e3",x"48",x"c3",x"ff"),
   393 => (x"50",x"c1",x"48",x"f5"),
   394 => (x"e8",x"87",x"0e",x"5e"),
   395 => (x"5b",x"5c",x"5d",x"0e"),
   396 => (x"1e",x"71",x"4a",x"c0"),
   397 => (x"4d",x"e3",x"48",x"c3"),
   398 => (x"ff",x"50",x"e7",x"48"),
   399 => (x"c2",x"50",x"eb",x"48"),
   400 => (x"c7",x"50",x"e3",x"48"),
   401 => (x"c3",x"ff",x"50",x"72"),
   402 => (x"1e",x"c0",x"ff",x"f0"),
   403 => (x"c1",x"d1",x"49",x"f2"),
   404 => (x"ce",x"87",x"c4",x"86"),
   405 => (x"70",x"98",x"05",x"c1"),
   406 => (x"c9",x"87",x"c5",x"ee"),
   407 => (x"cd",x"df",x"4b",x"e3"),
   408 => (x"48",x"c3",x"ff",x"50"),
   409 => (x"e3",x"97",x"bf",x"48"),
   410 => (x"c4",x"a6",x"58",x"6e"),
   411 => (x"49",x"c3",x"ff",x"99"),
   412 => (x"c3",x"fe",x"a9",x"05"),
   413 => (x"de",x"87",x"c0",x"4c"),
   414 => (x"ef",x"fd",x"87",x"d4"),
   415 => (x"66",x"08",x"78",x"08"),
   416 => (x"d4",x"66",x"48",x"c4"),
   417 => (x"80",x"d8",x"a6",x"58"),
   418 => (x"c1",x"84",x"c2",x"c0"),
   419 => (x"b7",x"ac",x"04",x"e7"),
   420 => (x"87",x"c1",x"4b",x"4d"),
   421 => (x"c1",x"8b",x"05",x"ff"),
   422 => (x"c5",x"87",x"e3",x"48"),
   423 => (x"c3",x"ff",x"50",x"e7"),
   424 => (x"48",x"c3",x"50",x"75"),
   425 => (x"48",x"26",x"f3",x"e5"),
   426 => (x"87",x"1e",x"73",x"1e"),
   427 => (x"71",x"4b",x"73",x"49"),
   428 => (x"d8",x"29",x"c3",x"ff"),
   429 => (x"99",x"73",x"4a",x"c8"),
   430 => (x"2a",x"cf",x"fc",x"c0"),
   431 => (x"9a",x"72",x"b1",x"73"),
   432 => (x"4a",x"c8",x"32",x"c0"),
   433 => (x"ff",x"f0",x"c0",x"c0"),
   434 => (x"9a",x"72",x"b1",x"73"),
   435 => (x"4a",x"d8",x"32",x"ff"),
   436 => (x"c0",x"c0",x"c0",x"c0"),
   437 => (x"9a",x"72",x"b1",x"71"),
   438 => (x"48",x"c4",x"87",x"26"),
   439 => (x"4d",x"26",x"4c",x"26"),
   440 => (x"4b",x"26",x"4f",x"1e"),
   441 => (x"73",x"1e",x"71",x"4b"),
   442 => (x"73",x"49",x"c8",x"29"),
   443 => (x"c3",x"ff",x"99",x"73"),
   444 => (x"4a",x"c8",x"32",x"cf"),
   445 => (x"fc",x"c0",x"9a",x"72"),
   446 => (x"b1",x"71",x"48",x"e2"),
   447 => (x"87",x"0e",x"5e",x"5b"),
   448 => (x"5c",x"0e",x"71",x"4b"),
   449 => (x"c0",x"4c",x"d0",x"66"),
   450 => (x"48",x"c0",x"b7",x"a8"),
   451 => (x"06",x"c0",x"e3",x"87"),
   452 => (x"13",x"4a",x"cc",x"66"),
   453 => (x"97",x"bf",x"49",x"cc"),
   454 => (x"66",x"48",x"c1",x"80"),
   455 => (x"d0",x"a6",x"58",x"71"),
   456 => (x"b7",x"aa",x"02",x"c4"),
   457 => (x"87",x"c1",x"48",x"cc"),
   458 => (x"87",x"c1",x"84",x"d0"),
   459 => (x"66",x"b7",x"ac",x"04"),
   460 => (x"ff",x"dd",x"87",x"c0"),
   461 => (x"48",x"c2",x"87",x"26"),
   462 => (x"4d",x"26",x"4c",x"26"),
   463 => (x"4b",x"26",x"4f",x"0e"),
   464 => (x"5e",x"5b",x"5c",x"0e"),
   465 => (x"1e",x"c1",x"ce",x"c2"),
   466 => (x"48",x"ff",x"78",x"c1"),
   467 => (x"cd",x"d2",x"48",x"c0"),
   468 => (x"78",x"c0",x"ea",x"e4"),
   469 => (x"49",x"da",x"cf",x"87"),
   470 => (x"c1",x"c5",x"ca",x"1e"),
   471 => (x"c0",x"49",x"fb",x"c9"),
   472 => (x"87",x"c4",x"86",x"70"),
   473 => (x"98",x"05",x"c5",x"87"),
   474 => (x"c0",x"48",x"ca",x"f0"),
   475 => (x"87",x"c0",x"4b",x"c1"),
   476 => (x"cd",x"fe",x"48",x"c1"),
   477 => (x"78",x"c8",x"1e",x"c0"),
   478 => (x"ea",x"f1",x"1e",x"c1"),
   479 => (x"c6",x"c0",x"49",x"fd"),
   480 => (x"fb",x"87",x"c8",x"86"),
   481 => (x"70",x"98",x"05",x"c6"),
   482 => (x"87",x"c1",x"cd",x"fe"),
   483 => (x"48",x"c0",x"78",x"c8"),
   484 => (x"1e",x"c0",x"ea",x"fa"),
   485 => (x"1e",x"c1",x"c6",x"dc"),
   486 => (x"49",x"fd",x"e1",x"87"),
   487 => (x"c8",x"86",x"70",x"98"),
   488 => (x"05",x"c6",x"87",x"c1"),
   489 => (x"cd",x"fe",x"48",x"c0"),
   490 => (x"78",x"c8",x"1e",x"c0"),
   491 => (x"eb",x"c3",x"1e",x"c1"),
   492 => (x"c6",x"dc",x"49",x"fd"),
   493 => (x"c7",x"87",x"c8",x"86"),
   494 => (x"70",x"98",x"05",x"c5"),
   495 => (x"87",x"c0",x"48",x"c9"),
   496 => (x"db",x"87",x"c1",x"cd"),
   497 => (x"fe",x"bf",x"1e",x"c0"),
   498 => (x"eb",x"cc",x"1e",x"c0"),
   499 => (x"e3",x"f5",x"87",x"c8"),
   500 => (x"86",x"c1",x"cd",x"fe"),
   501 => (x"bf",x"02",x"c1",x"ed"),
   502 => (x"87",x"c1",x"c5",x"ca"),
   503 => (x"4a",x"48",x"c6",x"fe"),
   504 => (x"a0",x"4c",x"c1",x"cc"),
   505 => (x"d0",x"bf",x"4b",x"c1"),
   506 => (x"cd",x"c8",x"9f",x"bf"),
   507 => (x"49",x"c4",x"a6",x"5a"),
   508 => (x"c5",x"d6",x"ea",x"a9"),
   509 => (x"05",x"c0",x"cc",x"87"),
   510 => (x"c8",x"a4",x"4a",x"6a"),
   511 => (x"49",x"fa",x"e9",x"87"),
   512 => (x"70",x"4b",x"db",x"87"),
   513 => (x"c7",x"fe",x"a2",x"49"),
   514 => (x"9f",x"69",x"49",x"ca"),
   515 => (x"e9",x"d5",x"a9",x"02"),
   516 => (x"c0",x"cc",x"87",x"c0"),
   517 => (x"e8",x"e1",x"49",x"d7"),
   518 => (x"cd",x"87",x"c0",x"48"),
   519 => (x"c7",x"fe",x"87",x"73"),
   520 => (x"1e",x"c0",x"e8",x"ff"),
   521 => (x"1e",x"c0",x"e2",x"db"),
   522 => (x"87",x"c1",x"c5",x"ca"),
   523 => (x"1e",x"73",x"49",x"f7"),
   524 => (x"f8",x"87",x"cc",x"86"),
   525 => (x"70",x"98",x"05",x"c0"),
   526 => (x"c5",x"87",x"c0",x"48"),
   527 => (x"c7",x"de",x"87",x"c0"),
   528 => (x"e9",x"d7",x"49",x"d6"),
   529 => (x"e1",x"87",x"c0",x"eb"),
   530 => (x"df",x"1e",x"c0",x"e1"),
   531 => (x"f6",x"87",x"c8",x"1e"),
   532 => (x"c0",x"eb",x"f7",x"1e"),
   533 => (x"c1",x"c6",x"dc",x"49"),
   534 => (x"fa",x"e2",x"87",x"cc"),
   535 => (x"86",x"70",x"98",x"05"),
   536 => (x"c0",x"c9",x"87",x"c1"),
   537 => (x"cd",x"d2",x"48",x"c1"),
   538 => (x"78",x"c0",x"e4",x"87"),
   539 => (x"c8",x"1e",x"c0",x"ec"),
   540 => (x"c0",x"1e",x"c1",x"c6"),
   541 => (x"c0",x"49",x"fa",x"c4"),
   542 => (x"87",x"c8",x"86",x"70"),
   543 => (x"98",x"02",x"c0",x"cf"),
   544 => (x"87",x"c0",x"e9",x"fe"),
   545 => (x"1e",x"c0",x"e0",x"fb"),
   546 => (x"87",x"c4",x"86",x"c0"),
   547 => (x"48",x"c6",x"cd",x"87"),
   548 => (x"c1",x"cd",x"c8",x"97"),
   549 => (x"bf",x"49",x"c1",x"d5"),
   550 => (x"a9",x"05",x"c0",x"cd"),
   551 => (x"87",x"c1",x"cd",x"c9"),
   552 => (x"97",x"bf",x"49",x"c2"),
   553 => (x"ea",x"a9",x"02",x"c0"),
   554 => (x"c5",x"87",x"c0",x"48"),
   555 => (x"c5",x"ee",x"87",x"c1"),
   556 => (x"c5",x"ca",x"97",x"bf"),
   557 => (x"49",x"c3",x"e9",x"a9"),
   558 => (x"02",x"c0",x"d2",x"87"),
   559 => (x"c1",x"c5",x"ca",x"97"),
   560 => (x"bf",x"49",x"c3",x"eb"),
   561 => (x"a9",x"02",x"c0",x"c5"),
   562 => (x"87",x"c0",x"48",x"c5"),
   563 => (x"cf",x"87",x"c1",x"c5"),
   564 => (x"d5",x"97",x"bf",x"49"),
   565 => (x"71",x"99",x"05",x"c0"),
   566 => (x"cc",x"87",x"c1",x"c5"),
   567 => (x"d6",x"97",x"bf",x"49"),
   568 => (x"c2",x"a9",x"02",x"c0"),
   569 => (x"c5",x"87",x"c0",x"48"),
   570 => (x"c4",x"f2",x"87",x"c1"),
   571 => (x"c5",x"d7",x"97",x"bf"),
   572 => (x"48",x"c1",x"cd",x"ce"),
   573 => (x"58",x"c1",x"cd",x"ca"),
   574 => (x"bf",x"48",x"c1",x"88"),
   575 => (x"c1",x"cd",x"d2",x"58"),
   576 => (x"c1",x"c5",x"d8",x"97"),
   577 => (x"bf",x"49",x"73",x"81"),
   578 => (x"c1",x"c5",x"d9",x"97"),
   579 => (x"bf",x"4a",x"c8",x"32"),
   580 => (x"c1",x"cd",x"de",x"48"),
   581 => (x"72",x"a1",x"78",x"c1"),
   582 => (x"c5",x"da",x"97",x"bf"),
   583 => (x"48",x"c1",x"cd",x"f6"),
   584 => (x"58",x"c1",x"cd",x"d2"),
   585 => (x"bf",x"02",x"c2",x"e2"),
   586 => (x"87",x"c8",x"1e",x"c0"),
   587 => (x"ea",x"db",x"1e",x"c1"),
   588 => (x"c6",x"dc",x"49",x"f7"),
   589 => (x"c7",x"87",x"c8",x"86"),
   590 => (x"70",x"98",x"02",x"c0"),
   591 => (x"c5",x"87",x"c0",x"48"),
   592 => (x"c3",x"da",x"87",x"c1"),
   593 => (x"cd",x"ca",x"bf",x"48"),
   594 => (x"c4",x"30",x"c1",x"cd"),
   595 => (x"fa",x"58",x"c1",x"cd"),
   596 => (x"ca",x"bf",x"4a",x"c1"),
   597 => (x"cd",x"f2",x"5a",x"c1"),
   598 => (x"c5",x"ef",x"97",x"bf"),
   599 => (x"49",x"c8",x"31",x"c1"),
   600 => (x"c5",x"ee",x"97",x"bf"),
   601 => (x"4b",x"73",x"a1",x"49"),
   602 => (x"c1",x"c5",x"f0",x"97"),
   603 => (x"bf",x"4b",x"d0",x"33"),
   604 => (x"73",x"a1",x"49",x"c1"),
   605 => (x"c5",x"f1",x"97",x"bf"),
   606 => (x"4b",x"d8",x"33",x"73"),
   607 => (x"a1",x"49",x"c1",x"cd"),
   608 => (x"fe",x"59",x"c1",x"cd"),
   609 => (x"f2",x"bf",x"91",x"c1"),
   610 => (x"cd",x"de",x"bf",x"81"),
   611 => (x"c1",x"cd",x"e6",x"59"),
   612 => (x"c1",x"c5",x"f7",x"97"),
   613 => (x"bf",x"4b",x"c8",x"33"),
   614 => (x"c1",x"c5",x"f6",x"97"),
   615 => (x"bf",x"4c",x"74",x"a3"),
   616 => (x"4b",x"c1",x"c5",x"f8"),
   617 => (x"97",x"bf",x"4c",x"d0"),
   618 => (x"34",x"74",x"a3",x"4b"),
   619 => (x"c1",x"c5",x"f9",x"97"),
   620 => (x"bf",x"4c",x"cf",x"9c"),
   621 => (x"d8",x"34",x"74",x"a3"),
   622 => (x"4b",x"c1",x"cd",x"ea"),
   623 => (x"5b",x"c2",x"8b",x"73"),
   624 => (x"92",x"c1",x"cd",x"ea"),
   625 => (x"48",x"72",x"a1",x"78"),
   626 => (x"c1",x"d0",x"87",x"c1"),
   627 => (x"c5",x"dc",x"97",x"bf"),
   628 => (x"49",x"c8",x"31",x"c1"),
   629 => (x"c5",x"db",x"97",x"bf"),
   630 => (x"4a",x"72",x"a1",x"49"),
   631 => (x"c1",x"cd",x"fa",x"59"),
   632 => (x"c5",x"31",x"c7",x"ff"),
   633 => (x"81",x"c9",x"29",x"c1"),
   634 => (x"cd",x"f2",x"59",x"c1"),
   635 => (x"c5",x"e1",x"97",x"bf"),
   636 => (x"4a",x"c8",x"32",x"c1"),
   637 => (x"c5",x"e0",x"97",x"bf"),
   638 => (x"4b",x"73",x"a2",x"4a"),
   639 => (x"c1",x"cd",x"fe",x"5a"),
   640 => (x"c1",x"cd",x"f2",x"bf"),
   641 => (x"92",x"c1",x"cd",x"de"),
   642 => (x"bf",x"82",x"c1",x"cd"),
   643 => (x"ee",x"5a",x"c1",x"cd"),
   644 => (x"e6",x"48",x"c0",x"78"),
   645 => (x"c1",x"cd",x"e2",x"48"),
   646 => (x"72",x"a1",x"78",x"c1"),
   647 => (x"48",x"26",x"f4",x"d8"),
   648 => (x"87",x"4e",x"6f",x"20"),
   649 => (x"70",x"61",x"72",x"74"),
   650 => (x"69",x"74",x"69",x"6f"),
   651 => (x"6e",x"20",x"73",x"69"),
   652 => (x"67",x"6e",x"61",x"74"),
   653 => (x"75",x"72",x"65",x"20"),
   654 => (x"66",x"6f",x"75",x"6e"),
   655 => (x"64",x"0a",x"00",x"52"),
   656 => (x"65",x"61",x"64",x"69"),
   657 => (x"6e",x"67",x"20",x"62"),
   658 => (x"6f",x"6f",x"74",x"20"),
   659 => (x"73",x"65",x"63",x"74"),
   660 => (x"6f",x"72",x"20",x"25"),
   661 => (x"64",x"0a",x"00",x"52"),
   662 => (x"65",x"61",x"64",x"20"),
   663 => (x"62",x"6f",x"6f",x"74"),
   664 => (x"20",x"73",x"65",x"63"),
   665 => (x"74",x"6f",x"72",x"20"),
   666 => (x"66",x"72",x"6f",x"6d"),
   667 => (x"20",x"66",x"69",x"72"),
   668 => (x"73",x"74",x"20",x"70"),
   669 => (x"61",x"72",x"74",x"69"),
   670 => (x"74",x"69",x"6f",x"6e"),
   671 => (x"0a",x"00",x"55",x"6e"),
   672 => (x"73",x"75",x"70",x"70"),
   673 => (x"6f",x"72",x"74",x"65"),
   674 => (x"64",x"20",x"70",x"61"),
   675 => (x"72",x"74",x"69",x"74"),
   676 => (x"69",x"6f",x"6e",x"20"),
   677 => (x"74",x"79",x"70",x"65"),
   678 => (x"21",x"0d",x"00",x"46"),
   679 => (x"41",x"54",x"33",x"32"),
   680 => (x"20",x"20",x"20",x"00"),
   681 => (x"52",x"65",x"61",x"64"),
   682 => (x"69",x"6e",x"67",x"20"),
   683 => (x"4d",x"42",x"52",x"0a"),
   684 => (x"00",x"46",x"41",x"54"),
   685 => (x"31",x"36",x"20",x"20"),
   686 => (x"20",x"00",x"46",x"41"),
   687 => (x"54",x"33",x"32",x"20"),
   688 => (x"20",x"20",x"00",x"46"),
   689 => (x"41",x"54",x"31",x"32"),
   690 => (x"20",x"20",x"20",x"00"),
   691 => (x"50",x"61",x"72",x"74"),
   692 => (x"69",x"74",x"69",x"6f"),
   693 => (x"6e",x"63",x"6f",x"75"),
   694 => (x"6e",x"74",x"20",x"25"),
   695 => (x"64",x"0a",x"00",x"48"),
   696 => (x"75",x"6e",x"74",x"69"),
   697 => (x"6e",x"67",x"20",x"66"),
   698 => (x"6f",x"72",x"20",x"66"),
   699 => (x"69",x"6c",x"65",x"73"),
   700 => (x"79",x"73",x"74",x"65"),
   701 => (x"6d",x"0a",x"00",x"46"),
   702 => (x"41",x"54",x"33",x"32"),
   703 => (x"20",x"20",x"20",x"00"),
   704 => (x"46",x"41",x"54",x"31"),
   705 => (x"36",x"20",x"20",x"20"),
   706 => (x"00",x"52",x"65",x"61"),
   707 => (x"64",x"69",x"6e",x"67"),
   708 => (x"20",x"64",x"69",x"72"),
   709 => (x"65",x"63",x"74",x"6f"),
   710 => (x"72",x"79",x"20",x"73"),
   711 => (x"65",x"63",x"74",x"6f"),
   712 => (x"72",x"20",x"25",x"64"),
   713 => (x"0a",x"00",x"66",x"69"),
   714 => (x"6c",x"65",x"20",x"22"),
   715 => (x"25",x"73",x"22",x"20"),
   716 => (x"66",x"6f",x"75",x"6e"),
   717 => (x"64",x"0d",x"00",x"47"),
   718 => (x"65",x"74",x"46",x"41"),
   719 => (x"54",x"4c",x"69",x"6e"),
   720 => (x"6b",x"20",x"72",x"65"),
   721 => (x"74",x"75",x"72",x"6e"),
   722 => (x"65",x"64",x"20",x"25"),
   723 => (x"64",x"0a",x"00",x"43"),
   724 => (x"61",x"6e",x"27",x"74"),
   725 => (x"20",x"6f",x"70",x"65"),
   726 => (x"6e",x"20",x"25",x"73"),
   727 => (x"0a",x"00",x"0e",x"5e"),
   728 => (x"5b",x"5c",x"5d",x"0e"),
   729 => (x"71",x"4a",x"c1",x"cd"),
   730 => (x"d2",x"bf",x"02",x"cc"),
   731 => (x"87",x"72",x"4b",x"c7"),
   732 => (x"b7",x"2b",x"72",x"4c"),
   733 => (x"c1",x"ff",x"9c",x"ca"),
   734 => (x"87",x"72",x"4b",x"c8"),
   735 => (x"b7",x"2b",x"72",x"4c"),
   736 => (x"c3",x"ff",x"9c",x"c1"),
   737 => (x"ce",x"c2",x"bf",x"ab"),
   738 => (x"02",x"de",x"87",x"c1"),
   739 => (x"c5",x"ca",x"1e",x"c1"),
   740 => (x"cd",x"de",x"bf",x"49"),
   741 => (x"73",x"81",x"ea",x"d1"),
   742 => (x"87",x"c4",x"86",x"70"),
   743 => (x"98",x"05",x"c5",x"87"),
   744 => (x"c0",x"48",x"c0",x"f6"),
   745 => (x"87",x"c1",x"ce",x"c6"),
   746 => (x"5b",x"c1",x"cd",x"d2"),
   747 => (x"bf",x"02",x"d9",x"87"),
   748 => (x"74",x"4a",x"c4",x"92"),
   749 => (x"c1",x"c5",x"ca",x"82"),
   750 => (x"6a",x"49",x"eb",x"ec"),
   751 => (x"87",x"70",x"49",x"71"),
   752 => (x"4d",x"cf",x"ff",x"ff"),
   753 => (x"ff",x"ff",x"9d",x"d0"),
   754 => (x"87",x"74",x"4a",x"c2"),
   755 => (x"92",x"c1",x"c5",x"ca"),
   756 => (x"82",x"9f",x"6a",x"49"),
   757 => (x"ec",x"cc",x"87",x"70"),
   758 => (x"4d",x"75",x"48",x"ed"),
   759 => (x"d9",x"87",x"0e",x"5e"),
   760 => (x"5b",x"5c",x"5d",x"0e"),
   761 => (x"f4",x"86",x"71",x"4c"),
   762 => (x"c0",x"4b",x"c1",x"ce"),
   763 => (x"c2",x"48",x"ff",x"78"),
   764 => (x"c1",x"cd",x"e6",x"bf"),
   765 => (x"4d",x"c1",x"cd",x"ea"),
   766 => (x"bf",x"7e",x"c1",x"cd"),
   767 => (x"d2",x"bf",x"02",x"c9"),
   768 => (x"87",x"c1",x"cd",x"ca"),
   769 => (x"bf",x"4a",x"c4",x"32"),
   770 => (x"c7",x"87",x"c1",x"cd"),
   771 => (x"ee",x"bf",x"4a",x"c4"),
   772 => (x"32",x"c8",x"a6",x"5a"),
   773 => (x"c8",x"a6",x"48",x"c0"),
   774 => (x"78",x"c4",x"66",x"48"),
   775 => (x"c0",x"a8",x"06",x"c3"),
   776 => (x"cf",x"87",x"c8",x"66"),
   777 => (x"49",x"cf",x"99",x"05"),
   778 => (x"c0",x"e3",x"87",x"6e"),
   779 => (x"1e",x"c0",x"ec",x"c9"),
   780 => (x"1e",x"d2",x"d0",x"87"),
   781 => (x"c1",x"c5",x"ca",x"1e"),
   782 => (x"cc",x"66",x"49",x"48"),
   783 => (x"c1",x"80",x"d0",x"a6"),
   784 => (x"58",x"71",x"49",x"e7"),
   785 => (x"e4",x"87",x"cc",x"86"),
   786 => (x"c1",x"c5",x"ca",x"4b"),
   787 => (x"c3",x"87",x"c0",x"e0"),
   788 => (x"83",x"97",x"6b",x"49"),
   789 => (x"71",x"99",x"02",x"c2"),
   790 => (x"c5",x"87",x"97",x"6b"),
   791 => (x"49",x"c3",x"e5",x"a9"),
   792 => (x"02",x"c1",x"fb",x"87"),
   793 => (x"cb",x"a3",x"49",x"97"),
   794 => (x"69",x"49",x"d8",x"99"),
   795 => (x"05",x"c1",x"ef",x"87"),
   796 => (x"cb",x"1e",x"c0",x"e0"),
   797 => (x"66",x"1e",x"73",x"49"),
   798 => (x"ea",x"c2",x"87",x"c8"),
   799 => (x"86",x"70",x"98",x"05"),
   800 => (x"c1",x"dc",x"87",x"dc"),
   801 => (x"a3",x"4a",x"6a",x"49"),
   802 => (x"e8",x"de",x"87",x"70"),
   803 => (x"4a",x"c4",x"a4",x"49"),
   804 => (x"72",x"79",x"da",x"a3"),
   805 => (x"4a",x"9f",x"6a",x"49"),
   806 => (x"e9",x"c8",x"87",x"c4"),
   807 => (x"a6",x"58",x"c1",x"cd"),
   808 => (x"d2",x"bf",x"02",x"d8"),
   809 => (x"87",x"d4",x"a3",x"4a"),
   810 => (x"9f",x"6a",x"49",x"e8"),
   811 => (x"f5",x"87",x"70",x"49"),
   812 => (x"c0",x"ff",x"ff",x"99"),
   813 => (x"71",x"48",x"d0",x"30"),
   814 => (x"c8",x"a6",x"58",x"c5"),
   815 => (x"87",x"c4",x"a6",x"48"),
   816 => (x"c0",x"78",x"c4",x"66"),
   817 => (x"4a",x"6e",x"82",x"c8"),
   818 => (x"a4",x"49",x"72",x"79"),
   819 => (x"c0",x"7c",x"dc",x"66"),
   820 => (x"1e",x"c0",x"ec",x"e6"),
   821 => (x"1e",x"cf",x"ec",x"87"),
   822 => (x"c8",x"86",x"c1",x"48"),
   823 => (x"c1",x"d0",x"87",x"c8"),
   824 => (x"66",x"48",x"c1",x"80"),
   825 => (x"cc",x"a6",x"58",x"c8"),
   826 => (x"66",x"48",x"c4",x"66"),
   827 => (x"a8",x"04",x"fc",x"f1"),
   828 => (x"87",x"c1",x"cd",x"d2"),
   829 => (x"bf",x"02",x"c0",x"f4"),
   830 => (x"87",x"75",x"49",x"f9"),
   831 => (x"e0",x"87",x"70",x"4d"),
   832 => (x"75",x"1e",x"c0",x"ec"),
   833 => (x"f7",x"1e",x"ce",x"fb"),
   834 => (x"87",x"c8",x"86",x"75"),
   835 => (x"49",x"cf",x"ff",x"ff"),
   836 => (x"ff",x"f8",x"99",x"a9"),
   837 => (x"02",x"d6",x"87",x"75"),
   838 => (x"49",x"c2",x"89",x"c1"),
   839 => (x"cd",x"ca",x"bf",x"91"),
   840 => (x"c1",x"cd",x"e2",x"bf"),
   841 => (x"48",x"71",x"80",x"c4"),
   842 => (x"a6",x"58",x"fb",x"e7"),
   843 => (x"87",x"c0",x"48",x"f4"),
   844 => (x"8e",x"e8",x"c3",x"87"),
   845 => (x"0e",x"5e",x"5b",x"5c"),
   846 => (x"5d",x"0e",x"1e",x"71"),
   847 => (x"4b",x"73",x"1e",x"c1"),
   848 => (x"ce",x"c6",x"49",x"fa"),
   849 => (x"d8",x"87",x"c4",x"86"),
   850 => (x"70",x"98",x"02",x"c1"),
   851 => (x"f7",x"87",x"c1",x"ce"),
   852 => (x"ca",x"bf",x"49",x"c7"),
   853 => (x"ff",x"81",x"c9",x"29"),
   854 => (x"c4",x"a6",x"59",x"c0"),
   855 => (x"4d",x"4c",x"6e",x"48"),
   856 => (x"c0",x"b7",x"a8",x"06"),
   857 => (x"c1",x"ed",x"87",x"c1"),
   858 => (x"cd",x"e2",x"bf",x"49"),
   859 => (x"c1",x"ce",x"ce",x"bf"),
   860 => (x"4a",x"c2",x"8a",x"c1"),
   861 => (x"cd",x"ca",x"bf",x"92"),
   862 => (x"72",x"a1",x"49",x"c1"),
   863 => (x"cd",x"ce",x"bf",x"4a"),
   864 => (x"74",x"9a",x"72",x"a1"),
   865 => (x"49",x"d4",x"66",x"1e"),
   866 => (x"71",x"49",x"e2",x"dd"),
   867 => (x"87",x"c4",x"86",x"70"),
   868 => (x"98",x"05",x"c5",x"87"),
   869 => (x"c0",x"48",x"c1",x"c0"),
   870 => (x"87",x"c1",x"84",x"c1"),
   871 => (x"cd",x"ce",x"bf",x"49"),
   872 => (x"74",x"99",x"05",x"cc"),
   873 => (x"87",x"c1",x"ce",x"ce"),
   874 => (x"bf",x"49",x"f6",x"f1"),
   875 => (x"87",x"c1",x"ce",x"d2"),
   876 => (x"58",x"d4",x"66",x"48"),
   877 => (x"c8",x"c0",x"80",x"d8"),
   878 => (x"a6",x"58",x"c1",x"85"),
   879 => (x"6e",x"b7",x"ad",x"04"),
   880 => (x"fe",x"e4",x"87",x"cf"),
   881 => (x"87",x"73",x"1e",x"c0"),
   882 => (x"ed",x"cf",x"1e",x"cb"),
   883 => (x"f6",x"87",x"c8",x"86"),
   884 => (x"c0",x"48",x"c5",x"87"),
   885 => (x"c1",x"ce",x"ca",x"bf"),
   886 => (x"48",x"26",x"e5",x"da"),
   887 => (x"87",x"1e",x"f3",x"09"),
   888 => (x"97",x"79",x"09",x"71"),
   889 => (x"48",x"26",x"4f",x"0e"),
   890 => (x"5e",x"5b",x"5c",x"0e"),
   891 => (x"71",x"4b",x"c0",x"4c"),
   892 => (x"13",x"4a",x"72",x"9a"),
   893 => (x"02",x"cd",x"87",x"72"),
   894 => (x"49",x"e2",x"87",x"c1"),
   895 => (x"84",x"13",x"4a",x"72"),
   896 => (x"9a",x"05",x"f3",x"87"),
   897 => (x"74",x"48",x"c2",x"87"),
   898 => (x"26",x"4d",x"26",x"4c"),
   899 => (x"26",x"4b",x"26",x"4f"),
   900 => (x"0e",x"5e",x"5b",x"5c"),
   901 => (x"5d",x"0e",x"fc",x"86"),
   902 => (x"71",x"4a",x"c0",x"e0"),
   903 => (x"66",x"4c",x"c1",x"ce"),
   904 => (x"d2",x"4b",x"c0",x"7e"),
   905 => (x"72",x"9a",x"05",x"ce"),
   906 => (x"87",x"c1",x"ce",x"d3"),
   907 => (x"4b",x"c1",x"ce",x"d2"),
   908 => (x"48",x"c0",x"f0",x"50"),
   909 => (x"c1",x"d2",x"87",x"72"),
   910 => (x"9a",x"02",x"c0",x"e9"),
   911 => (x"87",x"d4",x"66",x"4d"),
   912 => (x"72",x"1e",x"72",x"49"),
   913 => (x"75",x"4a",x"ca",x"cf"),
   914 => (x"87",x"26",x"4a",x"c0"),
   915 => (x"fa",x"fa",x"81",x"11"),
   916 => (x"53",x"71",x"1e",x"72"),
   917 => (x"49",x"75",x"4a",x"c9"),
   918 => (x"fe",x"87",x"70",x"4a"),
   919 => (x"26",x"49",x"c1",x"8c"),
   920 => (x"72",x"9a",x"05",x"ff"),
   921 => (x"da",x"87",x"c0",x"b7"),
   922 => (x"ac",x"06",x"dd",x"87"),
   923 => (x"c0",x"e4",x"66",x"02"),
   924 => (x"c5",x"87",x"c0",x"f0"),
   925 => (x"4a",x"c3",x"87",x"c0"),
   926 => (x"e0",x"4a",x"73",x"0a"),
   927 => (x"97",x"7a",x"0a",x"c1"),
   928 => (x"83",x"8c",x"c0",x"b7"),
   929 => (x"ac",x"01",x"ff",x"e3"),
   930 => (x"87",x"c1",x"ce",x"d2"),
   931 => (x"ab",x"02",x"de",x"87"),
   932 => (x"d8",x"66",x"4c",x"dc"),
   933 => (x"66",x"1e",x"c1",x"8b"),
   934 => (x"97",x"6b",x"49",x"74"),
   935 => (x"0f",x"c4",x"86",x"6e"),
   936 => (x"48",x"c1",x"80",x"c4"),
   937 => (x"a6",x"58",x"c1",x"ce"),
   938 => (x"d2",x"ab",x"05",x"ff"),
   939 => (x"e5",x"87",x"6e",x"48"),
   940 => (x"fc",x"8e",x"26",x"4d"),
   941 => (x"26",x"4c",x"26",x"4b"),
   942 => (x"26",x"4f",x"30",x"31"),
   943 => (x"32",x"33",x"34",x"35"),
   944 => (x"36",x"37",x"38",x"39"),
   945 => (x"41",x"42",x"43",x"44"),
   946 => (x"45",x"46",x"00",x"0e"),
   947 => (x"5e",x"5b",x"5c",x"5d"),
   948 => (x"0e",x"71",x"4b",x"ff"),
   949 => (x"4d",x"13",x"4c",x"74"),
   950 => (x"9c",x"02",x"d8",x"87"),
   951 => (x"c1",x"85",x"d4",x"66"),
   952 => (x"1e",x"74",x"49",x"d4"),
   953 => (x"66",x"0f",x"c4",x"86"),
   954 => (x"74",x"a8",x"05",x"c7"),
   955 => (x"87",x"13",x"4c",x"74"),
   956 => (x"9c",x"05",x"e8",x"87"),
   957 => (x"75",x"48",x"26",x"4d"),
   958 => (x"26",x"4c",x"26",x"4b"),
   959 => (x"26",x"4f",x"0e",x"5e"),
   960 => (x"5b",x"5c",x"5d",x"0e"),
   961 => (x"e8",x"86",x"c4",x"a6"),
   962 => (x"59",x"c0",x"e8",x"66"),
   963 => (x"4d",x"c0",x"4c",x"c8"),
   964 => (x"a6",x"48",x"c0",x"78"),
   965 => (x"6e",x"97",x"bf",x"4b"),
   966 => (x"6e",x"48",x"c1",x"80"),
   967 => (x"c4",x"a6",x"58",x"73"),
   968 => (x"9b",x"02",x"c6",x"d3"),
   969 => (x"87",x"c8",x"66",x"02"),
   970 => (x"c5",x"db",x"87",x"cc"),
   971 => (x"a6",x"48",x"c0",x"78"),
   972 => (x"fc",x"80",x"c0",x"78"),
   973 => (x"73",x"4a",x"c0",x"e0"),
   974 => (x"8a",x"02",x"c3",x"c6"),
   975 => (x"87",x"c3",x"8a",x"02"),
   976 => (x"c3",x"c0",x"87",x"c2"),
   977 => (x"8a",x"02",x"c2",x"e8"),
   978 => (x"87",x"c2",x"8a",x"02"),
   979 => (x"c2",x"f4",x"87",x"c4"),
   980 => (x"8a",x"02",x"c2",x"ee"),
   981 => (x"87",x"c2",x"8a",x"02"),
   982 => (x"c2",x"e8",x"87",x"c3"),
   983 => (x"8a",x"02",x"c2",x"ea"),
   984 => (x"87",x"d4",x"8a",x"02"),
   985 => (x"c0",x"f6",x"87",x"d4"),
   986 => (x"8a",x"02",x"c1",x"c0"),
   987 => (x"87",x"ca",x"8a",x"02"),
   988 => (x"c0",x"f2",x"87",x"c1"),
   989 => (x"8a",x"02",x"c1",x"e1"),
   990 => (x"87",x"c1",x"8a",x"02"),
   991 => (x"df",x"87",x"c8",x"8a"),
   992 => (x"02",x"c1",x"ce",x"87"),
   993 => (x"c4",x"8a",x"02",x"c0"),
   994 => (x"e3",x"87",x"c3",x"8a"),
   995 => (x"02",x"c0",x"e5",x"87"),
   996 => (x"c2",x"8a",x"02",x"c8"),
   997 => (x"87",x"c3",x"8a",x"02"),
   998 => (x"d3",x"87",x"c1",x"fa"),
   999 => (x"87",x"cc",x"a6",x"48"),
  1000 => (x"ca",x"78",x"c2",x"d2"),
  1001 => (x"87",x"cc",x"a6",x"48"),
  1002 => (x"c2",x"78",x"c2",x"ca"),
  1003 => (x"87",x"cc",x"a6",x"48"),
  1004 => (x"d0",x"78",x"c2",x"c2"),
  1005 => (x"87",x"c0",x"f0",x"66"),
  1006 => (x"1e",x"c0",x"f0",x"66"),
  1007 => (x"1e",x"c4",x"85",x"75"),
  1008 => (x"4a",x"c4",x"8a",x"6a"),
  1009 => (x"49",x"fc",x"c3",x"87"),
  1010 => (x"c8",x"86",x"70",x"49"),
  1011 => (x"71",x"a4",x"4c",x"c1"),
  1012 => (x"e5",x"87",x"c8",x"a6"),
  1013 => (x"48",x"c1",x"78",x"c1"),
  1014 => (x"dd",x"87",x"c0",x"f0"),
  1015 => (x"66",x"1e",x"c4",x"85"),
  1016 => (x"75",x"4a",x"c4",x"8a"),
  1017 => (x"6a",x"49",x"c0",x"f0"),
  1018 => (x"66",x"0f",x"c4",x"86"),
  1019 => (x"c1",x"84",x"c1",x"c6"),
  1020 => (x"87",x"c0",x"f0",x"66"),
  1021 => (x"1e",x"c0",x"e5",x"49"),
  1022 => (x"c0",x"f0",x"66",x"0f"),
  1023 => (x"c4",x"86",x"c1",x"84"),
  1024 => (x"c0",x"f4",x"87",x"c8"),
  1025 => (x"a6",x"48",x"c1",x"78"),
  1026 => (x"c0",x"ec",x"87",x"d0"),
  1027 => (x"a6",x"48",x"c1",x"78"),
  1028 => (x"f8",x"80",x"c1",x"78"),
  1029 => (x"c0",x"e0",x"87",x"c0"),
  1030 => (x"f0",x"ab",x"06",x"da"),
  1031 => (x"87",x"c0",x"f9",x"ab"),
  1032 => (x"03",x"d4",x"87",x"d4"),
  1033 => (x"66",x"49",x"ca",x"91"),
  1034 => (x"73",x"4a",x"c0",x"f0"),
  1035 => (x"8a",x"d4",x"a6",x"48"),
  1036 => (x"72",x"a1",x"78",x"f4"),
  1037 => (x"80",x"c1",x"78",x"cc"),
  1038 => (x"66",x"02",x"c1",x"ea"),
  1039 => (x"87",x"c4",x"85",x"75"),
  1040 => (x"49",x"c4",x"89",x"a6"),
  1041 => (x"48",x"69",x"78",x"c1"),
  1042 => (x"e4",x"ab",x"05",x"d8"),
  1043 => (x"87",x"c4",x"66",x"48"),
  1044 => (x"c0",x"b7",x"a8",x"03"),
  1045 => (x"cf",x"87",x"c0",x"ed"),
  1046 => (x"49",x"f6",x"c1",x"87"),
  1047 => (x"c4",x"66",x"48",x"c0"),
  1048 => (x"08",x"88",x"c8",x"a6"),
  1049 => (x"58",x"d0",x"66",x"1e"),
  1050 => (x"d8",x"66",x"1e",x"c0"),
  1051 => (x"f8",x"66",x"1e",x"c0"),
  1052 => (x"f8",x"66",x"1e",x"dc"),
  1053 => (x"66",x"1e",x"d8",x"66"),
  1054 => (x"49",x"f6",x"d4",x"87"),
  1055 => (x"d4",x"86",x"70",x"49"),
  1056 => (x"71",x"a4",x"4c",x"c0"),
  1057 => (x"e1",x"87",x"c0",x"e5"),
  1058 => (x"ab",x"05",x"cf",x"87"),
  1059 => (x"d0",x"a6",x"48",x"c0"),
  1060 => (x"78",x"c4",x"80",x"c0"),
  1061 => (x"78",x"f4",x"80",x"c1"),
  1062 => (x"78",x"cc",x"87",x"c0"),
  1063 => (x"f0",x"66",x"1e",x"73"),
  1064 => (x"49",x"c0",x"f0",x"66"),
  1065 => (x"0f",x"c4",x"86",x"6e"),
  1066 => (x"97",x"bf",x"4b",x"6e"),
  1067 => (x"48",x"c1",x"80",x"c4"),
  1068 => (x"a6",x"58",x"73",x"9b"),
  1069 => (x"05",x"f9",x"ed",x"87"),
  1070 => (x"74",x"48",x"e8",x"8e"),
  1071 => (x"26",x"4d",x"26",x"4c"),
  1072 => (x"26",x"4b",x"26",x"4f"),
  1073 => (x"1e",x"c0",x"1e",x"c0"),
  1074 => (x"f7",x"dd",x"1e",x"d0"),
  1075 => (x"a6",x"1e",x"d0",x"66"),
  1076 => (x"49",x"f8",x"ea",x"87"),
  1077 => (x"f4",x"8e",x"26",x"4f"),
  1078 => (x"1e",x"73",x"1e",x"72"),
  1079 => (x"9a",x"02",x"c0",x"e7"),
  1080 => (x"87",x"c0",x"48",x"c1"),
  1081 => (x"4b",x"72",x"a9",x"06"),
  1082 => (x"d1",x"87",x"72",x"82"),
  1083 => (x"06",x"c9",x"87",x"73"),
  1084 => (x"83",x"72",x"a9",x"01"),
  1085 => (x"f4",x"87",x"c3",x"87"),
  1086 => (x"c1",x"b2",x"3a",x"72"),
  1087 => (x"a9",x"03",x"89",x"73"),
  1088 => (x"80",x"07",x"c1",x"2a"),
  1089 => (x"2b",x"05",x"f3",x"87"),
  1090 => (x"26",x"4b",x"26",x"4f"),
  1091 => (x"1e",x"75",x"1e",x"c4"),
  1092 => (x"4d",x"71",x"b7",x"a1"),
  1093 => (x"04",x"ff",x"b9",x"c1"),
  1094 => (x"81",x"c3",x"bd",x"07"),
  1095 => (x"72",x"b7",x"a2",x"04"),
  1096 => (x"ff",x"ba",x"c1",x"82"),
  1097 => (x"c1",x"bd",x"07",x"fe"),
  1098 => (x"ee",x"87",x"c1",x"2d"),
  1099 => (x"04",x"ff",x"b8",x"c1"),
  1100 => (x"80",x"07",x"2d",x"04"),
  1101 => (x"ff",x"b9",x"c1",x"81"),
  1102 => (x"07",x"26",x"4d",x"26"),
  1103 => (x"4f",x"26",x"4d",x"26"),
	others => (others => x"00")
);

-- Xilinx XST attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "no_rw_check";

-- Altera Quartus attributes
attribute ramstyle: string;
attribute ramstyle of ram: signal is "no_rw_check";

signal q_local : word_t;

begin
    
	process(clk,q_local)
	begin

		q(31 downto 24)<=q_local(0);
		q(23 downto 16)<=q_local(1);
		q(15 downto 8)<=q_local(2);
		q(7 downto 0)<=q_local(3);

		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel(3) = '1') then
					ram(to_integer(unsigned(addr)))(3) <= d(7 downto 0);
				end if;
				if bytesel(2) = '1' then
					ram(to_integer(unsigned(addr)))(2) <= d(15 downto 8);
				end if;
				if bytesel(1) = '1' then
					ram(to_integer(unsigned(addr)))(1) <= d(23 downto 16);
				end if;
				if bytesel(0) = '1' then
					ram(to_integer(unsigned(addr)))(0) <= d(31 downto 24);
				end if;
			end if;
			q_local <= ram(to_integer(unsigned(addr)));
		end if;
	end process;

end arch;

