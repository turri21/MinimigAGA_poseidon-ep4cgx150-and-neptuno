library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM-2 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111";
	-- Second port
	addr2 : in std_logic_vector(maxAddrBitBRAM-2 downto 0) := (others=>'0');
	q2 : out std_logic_vector(31 downto 0);
	d2 : in std_logic_vector(31 downto 0) := X"00000000";
	we2 : in std_logic := '0';
	bytesel2 : in std_logic_vector(3 downto 0) := "1111"	
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
type ram_type is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

signal ram : ram_type :=
(
     0 => (x"01",x"da",x"87",x"04"),
     1 => (x"dd",x"87",x"0e",x"58"),
     2 => (x"5e",x"59",x"5a",x"0e"),
     3 => (x"27",x"00",x"00",x"00"),
     4 => (x"2c",x"0f",x"26",x"4a"),
     5 => (x"26",x"49",x"26",x"48"),
     6 => (x"ff",x"80",x"26",x"08"),
     7 => (x"4f",x"27",x"00",x"00"),
     8 => (x"00",x"2d",x"4f",x"27"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"4f",x"00",x"fd",x"87"),
    11 => (x"4f",x"c1",x"cd",x"e0"),
    12 => (x"4e",x"c9",x"c0",x"86"),
    13 => (x"c1",x"cd",x"e0",x"49"),
    14 => (x"c1",x"c3",x"fc",x"48"),
    15 => (x"89",x"d0",x"89",x"03"),
    16 => (x"c0",x"40",x"40",x"40"),
    17 => (x"40",x"f6",x"87",x"d0"),
    18 => (x"81",x"05",x"c0",x"50"),
    19 => (x"c1",x"89",x"05",x"f9"),
    20 => (x"87",x"c1",x"c3",x"f9"),
    21 => (x"4d",x"c1",x"c3",x"f9"),
    22 => (x"4c",x"74",x"ad",x"02"),
    23 => (x"c4",x"87",x"24",x"0f"),
    24 => (x"f7",x"87",x"c2",x"df"),
    25 => (x"87",x"c1",x"c3",x"f9"),
    26 => (x"4d",x"c1",x"c3",x"f9"),
    27 => (x"4c",x"74",x"ad",x"02"),
    28 => (x"c6",x"87",x"c4",x"8c"),
    29 => (x"6c",x"0f",x"f5",x"87"),
    30 => (x"00",x"fd",x"87",x"0e"),
    31 => (x"5e",x"5b",x"5c",x"0e"),
    32 => (x"c4",x"c0",x"c0",x"c0"),
    33 => (x"4b",x"c9",x"c3",x"4c"),
    34 => (x"c9",x"d5",x"bf",x"4a"),
    35 => (x"49",x"c1",x"8a",x"71"),
    36 => (x"99",x"02",x"cf",x"87"),
    37 => (x"74",x"49",x"c1",x"84"),
    38 => (x"11",x"53",x"72",x"49"),
    39 => (x"c1",x"8a",x"71",x"99"),
    40 => (x"05",x"f1",x"87",x"c2"),
    41 => (x"87",x"26",x"4d",x"26"),
    42 => (x"4c",x"26",x"4b",x"26"),
    43 => (x"4f",x"1e",x"73",x"1e"),
    44 => (x"71",x"4b",x"e7",x"48"),
    45 => (x"c0",x"e0",x"50",x"e3"),
    46 => (x"48",x"c8",x"50",x"e3"),
    47 => (x"48",x"c6",x"50",x"e7"),
    48 => (x"48",x"c0",x"e1",x"50"),
    49 => (x"73",x"4a",x"c8",x"b7"),
    50 => (x"2a",x"c4",x"c0",x"c0"),
    51 => (x"c0",x"49",x"ca",x"81"),
    52 => (x"71",x"0a",x"97",x"7a"),
    53 => (x"73",x"4a",x"c3",x"ff"),
    54 => (x"9a",x"c4",x"c0",x"c0"),
    55 => (x"c0",x"49",x"cb",x"81"),
    56 => (x"71",x"0a",x"97",x"7a"),
    57 => (x"e7",x"48",x"c0",x"e0"),
    58 => (x"50",x"e3",x"48",x"c8"),
    59 => (x"50",x"e3",x"48",x"c0"),
    60 => (x"50",x"e7",x"48",x"c0"),
    61 => (x"e1",x"50",x"fe",x"f0"),
    62 => (x"87",x"1e",x"73",x"1e"),
    63 => (x"c2",x"c0",x"c0",x"4b"),
    64 => (x"0f",x"fe",x"e5",x"87"),
    65 => (x"1e",x"73",x"1e",x"eb"),
    66 => (x"48",x"c3",x"ef",x"50"),
    67 => (x"e7",x"48",x"c0",x"e0"),
    68 => (x"50",x"e3",x"48",x"c8"),
    69 => (x"50",x"e3",x"48",x"c6"),
    70 => (x"50",x"e7",x"48",x"c0"),
    71 => (x"e1",x"50",x"ff",x"c2"),
    72 => (x"48",x"c1",x"9f",x"78"),
    73 => (x"e7",x"48",x"c0",x"e0"),
    74 => (x"50",x"e3",x"48",x"c4"),
    75 => (x"50",x"e3",x"48",x"c2"),
    76 => (x"50",x"e7",x"48",x"c0"),
    77 => (x"e1",x"50",x"e7",x"48"),
    78 => (x"c0",x"e0",x"50",x"e3"),
    79 => (x"48",x"c8",x"50",x"e3"),
    80 => (x"48",x"c7",x"50",x"e7"),
    81 => (x"48",x"c0",x"e1",x"50"),
    82 => (x"fc",x"f0",x"87",x"c0"),
    83 => (x"ff",x"ff",x"49",x"fd"),
    84 => (x"db",x"87",x"c0",x"fc"),
    85 => (x"c0",x"4b",x"c8",x"cf"),
    86 => (x"49",x"c0",x"f1",x"c8"),
    87 => (x"87",x"d0",x"eb",x"87"),
    88 => (x"70",x"98",x"02",x"c1"),
    89 => (x"c3",x"87",x"c0",x"ff"),
    90 => (x"f0",x"4b",x"c7",x"f8"),
    91 => (x"49",x"c0",x"f0",x"f4"),
    92 => (x"87",x"d6",x"d9",x"87"),
    93 => (x"70",x"98",x"02",x"c0"),
    94 => (x"e6",x"87",x"c3",x"f0"),
    95 => (x"4b",x"c2",x"c0",x"c0"),
    96 => (x"1e",x"c6",x"fb",x"49"),
    97 => (x"c0",x"ed",x"ec",x"87"),
    98 => (x"c4",x"86",x"70",x"98"),
    99 => (x"02",x"c8",x"87",x"c3"),
   100 => (x"ff",x"4b",x"fd",x"e4"),
   101 => (x"87",x"d9",x"87",x"c7"),
   102 => (x"c7",x"49",x"c0",x"f0"),
   103 => (x"c7",x"87",x"d0",x"87"),
   104 => (x"c7",x"dc",x"49",x"c0"),
   105 => (x"ef",x"fe",x"87",x"c7"),
   106 => (x"87",x"c8",x"e5",x"49"),
   107 => (x"c0",x"ef",x"f5",x"87"),
   108 => (x"73",x"49",x"fb",x"f8"),
   109 => (x"87",x"fe",x"da",x"87"),
   110 => (x"fb",x"ee",x"87",x"38"),
   111 => (x"33",x"32",x"4f",x"53"),
   112 => (x"44",x"41",x"44",x"42"),
   113 => (x"49",x"4e",x"00",x"43"),
   114 => (x"61",x"6e",x"27",x"74"),
   115 => (x"20",x"6c",x"6f",x"61"),
   116 => (x"64",x"20",x"66",x"69"),
   117 => (x"72",x"6d",x"77",x"61"),
   118 => (x"72",x"65",x"0a",x"00"),
   119 => (x"55",x"6e",x"61",x"62"),
   120 => (x"6c",x"65",x"20",x"74"),
   121 => (x"6f",x"20",x"6c",x"6f"),
   122 => (x"63",x"61",x"74",x"65"),
   123 => (x"20",x"70",x"61",x"72"),
   124 => (x"74",x"69",x"74",x"69"),
   125 => (x"6f",x"6e",x"0a",x"00"),
   126 => (x"48",x"75",x"6e",x"74"),
   127 => (x"69",x"6e",x"67",x"20"),
   128 => (x"66",x"6f",x"72",x"20"),
   129 => (x"70",x"61",x"72",x"74"),
   130 => (x"69",x"74",x"69",x"6f"),
   131 => (x"6e",x"0a",x"00",x"49"),
   132 => (x"6e",x"69",x"74",x"69"),
   133 => (x"61",x"6c",x"69",x"7a"),
   134 => (x"69",x"6e",x"67",x"20"),
   135 => (x"53",x"44",x"20",x"63"),
   136 => (x"61",x"72",x"64",x"0a"),
   137 => (x"00",x"46",x"61",x"69"),
   138 => (x"6c",x"65",x"64",x"20"),
   139 => (x"74",x"6f",x"20",x"69"),
   140 => (x"6e",x"69",x"74",x"69"),
   141 => (x"61",x"6c",x"69",x"7a"),
   142 => (x"65",x"20",x"53",x"44"),
   143 => (x"20",x"63",x"61",x"72"),
   144 => (x"64",x"0a",x"00",x"00"),
   145 => (x"00",x"00",x"00",x"00"),
   146 => (x"00",x"00",x"08",x"33"),
   147 => (x"fc",x"0f",x"ff",x"00"),
   148 => (x"df",x"f1",x"80",x"60"),
   149 => (x"f6",x"00",x"00",x"00"),
   150 => (x"12",x"1e",x"e4",x"86"),
   151 => (x"e3",x"48",x"c3",x"ff"),
   152 => (x"50",x"e3",x"97",x"bf"),
   153 => (x"48",x"c4",x"a6",x"58"),
   154 => (x"70",x"49",x"c3",x"ff"),
   155 => (x"99",x"e3",x"48",x"c3"),
   156 => (x"ff",x"50",x"c8",x"31"),
   157 => (x"e3",x"97",x"bf",x"48"),
   158 => (x"c8",x"a6",x"58",x"c3"),
   159 => (x"ff",x"98",x"cc",x"a6"),
   160 => (x"58",x"70",x"b1",x"e3"),
   161 => (x"48",x"c3",x"ff",x"50"),
   162 => (x"c8",x"31",x"e3",x"97"),
   163 => (x"bf",x"48",x"d0",x"a6"),
   164 => (x"58",x"c3",x"ff",x"98"),
   165 => (x"d4",x"a6",x"58",x"70"),
   166 => (x"b1",x"e3",x"48",x"c3"),
   167 => (x"ff",x"50",x"c8",x"31"),
   168 => (x"e3",x"97",x"bf",x"48"),
   169 => (x"d8",x"a6",x"58",x"c3"),
   170 => (x"ff",x"98",x"dc",x"a6"),
   171 => (x"58",x"70",x"b1",x"71"),
   172 => (x"48",x"e4",x"8e",x"26"),
   173 => (x"4f",x"0e",x"5e",x"5b"),
   174 => (x"5c",x"0e",x"1e",x"71"),
   175 => (x"4a",x"49",x"c3",x"ff"),
   176 => (x"99",x"e3",x"09",x"97"),
   177 => (x"79",x"09",x"c1",x"c3"),
   178 => (x"fc",x"bf",x"05",x"c8"),
   179 => (x"87",x"d0",x"66",x"48"),
   180 => (x"c9",x"30",x"d4",x"a6"),
   181 => (x"58",x"d0",x"66",x"49"),
   182 => (x"d8",x"29",x"c3",x"ff"),
   183 => (x"99",x"e3",x"09",x"97"),
   184 => (x"79",x"09",x"d0",x"66"),
   185 => (x"49",x"d0",x"29",x"c3"),
   186 => (x"ff",x"99",x"e3",x"09"),
   187 => (x"97",x"79",x"09",x"d0"),
   188 => (x"66",x"49",x"c8",x"29"),
   189 => (x"c3",x"ff",x"99",x"e3"),
   190 => (x"09",x"97",x"79",x"09"),
   191 => (x"d0",x"66",x"49",x"c3"),
   192 => (x"ff",x"99",x"e3",x"09"),
   193 => (x"97",x"79",x"09",x"72"),
   194 => (x"49",x"d0",x"29",x"c3"),
   195 => (x"ff",x"99",x"e3",x"09"),
   196 => (x"97",x"79",x"09",x"97"),
   197 => (x"bf",x"48",x"c4",x"a6"),
   198 => (x"58",x"70",x"4b",x"c3"),
   199 => (x"ff",x"9b",x"c9",x"f0"),
   200 => (x"ff",x"4c",x"c3",x"ff"),
   201 => (x"ab",x"05",x"dc",x"87"),
   202 => (x"e3",x"48",x"c3",x"ff"),
   203 => (x"50",x"e3",x"97",x"bf"),
   204 => (x"48",x"c4",x"a6",x"58"),
   205 => (x"70",x"4b",x"c3",x"ff"),
   206 => (x"9b",x"c1",x"8c",x"02"),
   207 => (x"c6",x"87",x"c3",x"ff"),
   208 => (x"ab",x"02",x"e4",x"87"),
   209 => (x"73",x"4a",x"c4",x"b7"),
   210 => (x"2a",x"c0",x"f0",x"a2"),
   211 => (x"49",x"c0",x"e9",x"ca"),
   212 => (x"87",x"73",x"4a",x"cf"),
   213 => (x"9a",x"c0",x"f0",x"a2"),
   214 => (x"49",x"c0",x"e8",x"fe"),
   215 => (x"87",x"73",x"48",x"26"),
   216 => (x"c2",x"87",x"26",x"4d"),
   217 => (x"26",x"4c",x"26",x"4b"),
   218 => (x"26",x"4f",x"1e",x"c0"),
   219 => (x"49",x"e3",x"48",x"c3"),
   220 => (x"ff",x"50",x"c1",x"81"),
   221 => (x"c3",x"c8",x"b7",x"a9"),
   222 => (x"04",x"f2",x"87",x"26"),
   223 => (x"4f",x"1e",x"73",x"1e"),
   224 => (x"e8",x"87",x"c4",x"f8"),
   225 => (x"df",x"4b",x"c0",x"1e"),
   226 => (x"c0",x"ff",x"f0",x"c1"),
   227 => (x"f7",x"49",x"fc",x"e4"),
   228 => (x"87",x"c4",x"86",x"c1"),
   229 => (x"a8",x"05",x"c0",x"e8"),
   230 => (x"87",x"e3",x"48",x"c3"),
   231 => (x"ff",x"50",x"c1",x"c0"),
   232 => (x"c0",x"c0",x"c0",x"c0"),
   233 => (x"1e",x"c0",x"e1",x"f0"),
   234 => (x"c1",x"e9",x"49",x"fc"),
   235 => (x"c7",x"87",x"c4",x"86"),
   236 => (x"70",x"98",x"05",x"c9"),
   237 => (x"87",x"e3",x"48",x"c3"),
   238 => (x"ff",x"50",x"c1",x"48"),
   239 => (x"cb",x"87",x"fe",x"e9"),
   240 => (x"87",x"c1",x"8b",x"05"),
   241 => (x"fe",x"ff",x"87",x"c0"),
   242 => (x"48",x"fe",x"da",x"87"),
   243 => (x"43",x"4d",x"44",x"34"),
   244 => (x"31",x"20",x"25",x"64"),
   245 => (x"0a",x"00",x"43",x"4d"),
   246 => (x"44",x"35",x"35",x"20"),
   247 => (x"25",x"64",x"0a",x"00"),
   248 => (x"43",x"4d",x"44",x"34"),
   249 => (x"31",x"20",x"25",x"64"),
   250 => (x"0a",x"00",x"43",x"4d"),
   251 => (x"44",x"35",x"35",x"20"),
   252 => (x"25",x"64",x"0a",x"00"),
   253 => (x"69",x"6e",x"69",x"74"),
   254 => (x"20",x"25",x"64",x"0a"),
   255 => (x"20",x"20",x"00",x"69"),
   256 => (x"6e",x"69",x"74",x"20"),
   257 => (x"25",x"64",x"0a",x"20"),
   258 => (x"20",x"00",x"43",x"6d"),
   259 => (x"64",x"5f",x"69",x"6e"),
   260 => (x"69",x"74",x"0a",x"00"),
   261 => (x"43",x"4d",x"44",x"38"),
   262 => (x"5f",x"34",x"20",x"72"),
   263 => (x"65",x"73",x"70",x"6f"),
   264 => (x"6e",x"73",x"65",x"3a"),
   265 => (x"20",x"25",x"64",x"0a"),
   266 => (x"00",x"43",x"4d",x"44"),
   267 => (x"35",x"38",x"20",x"25"),
   268 => (x"64",x"0a",x"20",x"20"),
   269 => (x"00",x"43",x"4d",x"44"),
   270 => (x"35",x"38",x"5f",x"32"),
   271 => (x"20",x"25",x"64",x"0a"),
   272 => (x"20",x"20",x"00",x"43"),
   273 => (x"4d",x"44",x"35",x"38"),
   274 => (x"20",x"25",x"64",x"0a"),
   275 => (x"20",x"20",x"00",x"53"),
   276 => (x"44",x"48",x"43",x"20"),
   277 => (x"49",x"6e",x"69",x"74"),
   278 => (x"69",x"61",x"6c",x"69"),
   279 => (x"7a",x"61",x"74",x"69"),
   280 => (x"6f",x"6e",x"20",x"65"),
   281 => (x"72",x"72",x"6f",x"72"),
   282 => (x"21",x"0a",x"00",x"63"),
   283 => (x"6d",x"64",x"5f",x"43"),
   284 => (x"4d",x"44",x"38",x"20"),
   285 => (x"72",x"65",x"73",x"70"),
   286 => (x"6f",x"6e",x"73",x"65"),
   287 => (x"3a",x"20",x"25",x"64"),
   288 => (x"0a",x"00",x"52",x"65"),
   289 => (x"61",x"64",x"20",x"63"),
   290 => (x"6f",x"6d",x"6d",x"61"),
   291 => (x"6e",x"64",x"20",x"66"),
   292 => (x"61",x"69",x"6c",x"65"),
   293 => (x"64",x"20",x"61",x"74"),
   294 => (x"20",x"25",x"64",x"20"),
   295 => (x"28",x"25",x"64",x"29"),
   296 => (x"0a",x"00",x"1e",x"73"),
   297 => (x"1e",x"e3",x"48",x"c3"),
   298 => (x"ff",x"50",x"d0",x"ca"),
   299 => (x"49",x"c0",x"e3",x"f4"),
   300 => (x"87",x"d3",x"4b",x"c0"),
   301 => (x"1e",x"c0",x"ff",x"f0"),
   302 => (x"c1",x"c1",x"49",x"f7"),
   303 => (x"f7",x"87",x"c4",x"86"),
   304 => (x"70",x"98",x"05",x"c9"),
   305 => (x"87",x"e3",x"48",x"c3"),
   306 => (x"ff",x"50",x"c1",x"48"),
   307 => (x"cb",x"87",x"fa",x"d9"),
   308 => (x"87",x"c1",x"8b",x"05"),
   309 => (x"ff",x"dc",x"87",x"c0"),
   310 => (x"48",x"fa",x"ca",x"87"),
   311 => (x"1e",x"73",x"1e",x"1e"),
   312 => (x"fa",x"c7",x"87",x"c6"),
   313 => (x"ea",x"1e",x"c0",x"e1"),
   314 => (x"f0",x"c1",x"c8",x"49"),
   315 => (x"f7",x"c6",x"87",x"70"),
   316 => (x"4b",x"1e",x"d1",x"eb"),
   317 => (x"1e",x"c0",x"ee",x"c7"),
   318 => (x"87",x"cc",x"86",x"c1"),
   319 => (x"ab",x"02",x"c8",x"87"),
   320 => (x"fe",x"df",x"87",x"c0"),
   321 => (x"48",x"c1",x"ff",x"87"),
   322 => (x"f5",x"ce",x"87",x"70"),
   323 => (x"49",x"cf",x"ff",x"ff"),
   324 => (x"99",x"c6",x"ea",x"a9"),
   325 => (x"02",x"c8",x"87",x"fe"),
   326 => (x"c8",x"87",x"c0",x"48"),
   327 => (x"c1",x"e8",x"87",x"e3"),
   328 => (x"48",x"c3",x"ff",x"50"),
   329 => (x"c0",x"f1",x"4b",x"f9"),
   330 => (x"d3",x"87",x"70",x"98"),
   331 => (x"02",x"c1",x"c6",x"87"),
   332 => (x"c0",x"1e",x"c0",x"ff"),
   333 => (x"f0",x"c1",x"fa",x"49"),
   334 => (x"f5",x"fa",x"87",x"c4"),
   335 => (x"86",x"70",x"98",x"05"),
   336 => (x"c0",x"f3",x"87",x"e3"),
   337 => (x"48",x"c3",x"ff",x"50"),
   338 => (x"e3",x"97",x"bf",x"48"),
   339 => (x"c4",x"a6",x"58",x"70"),
   340 => (x"49",x"c3",x"ff",x"99"),
   341 => (x"e3",x"48",x"c3",x"ff"),
   342 => (x"50",x"e3",x"48",x"c3"),
   343 => (x"ff",x"50",x"e3",x"48"),
   344 => (x"c3",x"ff",x"50",x"e3"),
   345 => (x"48",x"c3",x"ff",x"50"),
   346 => (x"c1",x"c0",x"99",x"02"),
   347 => (x"c4",x"87",x"c1",x"48"),
   348 => (x"d5",x"87",x"c0",x"48"),
   349 => (x"d1",x"87",x"c2",x"ab"),
   350 => (x"05",x"c4",x"87",x"c0"),
   351 => (x"48",x"c8",x"87",x"c1"),
   352 => (x"8b",x"05",x"fe",x"e2"),
   353 => (x"87",x"c0",x"48",x"26"),
   354 => (x"f7",x"db",x"87",x"1e"),
   355 => (x"73",x"1e",x"c1",x"c3"),
   356 => (x"fc",x"48",x"c1",x"78"),
   357 => (x"eb",x"48",x"c3",x"ef"),
   358 => (x"50",x"c7",x"4b",x"e7"),
   359 => (x"48",x"c3",x"50",x"f7"),
   360 => (x"c8",x"87",x"e7",x"48"),
   361 => (x"c2",x"50",x"e3",x"48"),
   362 => (x"c3",x"ff",x"50",x"c0"),
   363 => (x"1e",x"c0",x"e5",x"d0"),
   364 => (x"c1",x"c0",x"49",x"f3"),
   365 => (x"ff",x"87",x"c4",x"86"),
   366 => (x"c1",x"a8",x"05",x"c1"),
   367 => (x"87",x"4b",x"c2",x"ab"),
   368 => (x"05",x"c5",x"87",x"c0"),
   369 => (x"48",x"c0",x"ef",x"87"),
   370 => (x"c1",x"8b",x"05",x"ff"),
   371 => (x"cd",x"87",x"fc",x"cb"),
   372 => (x"87",x"c1",x"c4",x"c0"),
   373 => (x"58",x"70",x"98",x"05"),
   374 => (x"cd",x"87",x"c1",x"1e"),
   375 => (x"c0",x"ff",x"f0",x"c1"),
   376 => (x"d0",x"49",x"f3",x"d0"),
   377 => (x"87",x"c4",x"86",x"e3"),
   378 => (x"48",x"c3",x"ff",x"50"),
   379 => (x"e7",x"48",x"c3",x"50"),
   380 => (x"e3",x"48",x"c3",x"ff"),
   381 => (x"50",x"c1",x"48",x"f5"),
   382 => (x"ec",x"87",x"0e",x"5e"),
   383 => (x"5b",x"5c",x"5d",x"0e"),
   384 => (x"1e",x"71",x"4a",x"c0"),
   385 => (x"4d",x"e3",x"48",x"c3"),
   386 => (x"ff",x"50",x"e7",x"48"),
   387 => (x"c2",x"50",x"eb",x"48"),
   388 => (x"c7",x"50",x"e3",x"48"),
   389 => (x"c3",x"ff",x"50",x"72"),
   390 => (x"1e",x"c0",x"ff",x"f0"),
   391 => (x"c1",x"d1",x"49",x"f2"),
   392 => (x"d3",x"87",x"c4",x"86"),
   393 => (x"70",x"98",x"05",x"c1"),
   394 => (x"c9",x"87",x"c5",x"ee"),
   395 => (x"cd",x"df",x"4b",x"e3"),
   396 => (x"48",x"c3",x"ff",x"50"),
   397 => (x"e3",x"97",x"bf",x"48"),
   398 => (x"c4",x"a6",x"58",x"70"),
   399 => (x"49",x"c3",x"ff",x"99"),
   400 => (x"c3",x"fe",x"a9",x"05"),
   401 => (x"de",x"87",x"c0",x"4c"),
   402 => (x"f0",x"ce",x"87",x"d4"),
   403 => (x"66",x"08",x"78",x"08"),
   404 => (x"d4",x"66",x"48",x"c4"),
   405 => (x"80",x"d8",x"a6",x"58"),
   406 => (x"c1",x"84",x"c2",x"c0"),
   407 => (x"b7",x"ac",x"04",x"e7"),
   408 => (x"87",x"c1",x"4b",x"4d"),
   409 => (x"c1",x"8b",x"05",x"ff"),
   410 => (x"c5",x"87",x"e3",x"48"),
   411 => (x"c3",x"ff",x"50",x"e7"),
   412 => (x"48",x"c3",x"50",x"75"),
   413 => (x"48",x"26",x"f3",x"e9"),
   414 => (x"87",x"1e",x"73",x"1e"),
   415 => (x"71",x"4b",x"49",x"d8"),
   416 => (x"29",x"c3",x"ff",x"99"),
   417 => (x"73",x"4a",x"c8",x"2a"),
   418 => (x"cf",x"fc",x"c0",x"9a"),
   419 => (x"72",x"b1",x"73",x"4a"),
   420 => (x"c8",x"32",x"c0",x"ff"),
   421 => (x"f0",x"c0",x"c0",x"9a"),
   422 => (x"72",x"b1",x"73",x"4a"),
   423 => (x"d8",x"32",x"ff",x"c0"),
   424 => (x"c0",x"c0",x"c0",x"9a"),
   425 => (x"72",x"b1",x"71",x"48"),
   426 => (x"c4",x"87",x"26",x"4d"),
   427 => (x"26",x"4c",x"26",x"4b"),
   428 => (x"26",x"4f",x"1e",x"73"),
   429 => (x"1e",x"71",x"4b",x"49"),
   430 => (x"c8",x"29",x"c3",x"ff"),
   431 => (x"99",x"73",x"4a",x"c8"),
   432 => (x"32",x"cf",x"fc",x"c0"),
   433 => (x"9a",x"72",x"b1",x"71"),
   434 => (x"48",x"e3",x"87",x"0e"),
   435 => (x"5e",x"5b",x"5c",x"0e"),
   436 => (x"71",x"4b",x"c0",x"4c"),
   437 => (x"d0",x"66",x"48",x"c0"),
   438 => (x"b7",x"a8",x"06",x"c0"),
   439 => (x"e3",x"87",x"13",x"4a"),
   440 => (x"cc",x"66",x"97",x"bf"),
   441 => (x"49",x"cc",x"66",x"48"),
   442 => (x"c1",x"80",x"d0",x"a6"),
   443 => (x"58",x"71",x"b7",x"aa"),
   444 => (x"02",x"c4",x"87",x"c1"),
   445 => (x"48",x"cc",x"87",x"c1"),
   446 => (x"84",x"d0",x"66",x"b7"),
   447 => (x"ac",x"04",x"ff",x"dd"),
   448 => (x"87",x"c0",x"48",x"c2"),
   449 => (x"87",x"26",x"4d",x"26"),
   450 => (x"4c",x"26",x"4b",x"26"),
   451 => (x"4f",x"0e",x"5e",x"5b"),
   452 => (x"5c",x"0e",x"1e",x"c1"),
   453 => (x"cc",x"fe",x"48",x"ff"),
   454 => (x"78",x"c1",x"cc",x"ce"),
   455 => (x"48",x"c0",x"78",x"c0"),
   456 => (x"e9",x"e8",x"49",x"d9"),
   457 => (x"ff",x"87",x"c1",x"c4"),
   458 => (x"c6",x"1e",x"c0",x"49"),
   459 => (x"fb",x"cb",x"87",x"c4"),
   460 => (x"86",x"70",x"98",x"05"),
   461 => (x"c5",x"87",x"c0",x"48"),
   462 => (x"ca",x"e6",x"87",x"c0"),
   463 => (x"4b",x"c1",x"cc",x"fa"),
   464 => (x"48",x"c1",x"78",x"c8"),
   465 => (x"1e",x"c0",x"e9",x"f5"),
   466 => (x"1e",x"c1",x"c4",x"fc"),
   467 => (x"49",x"fd",x"fb",x"87"),
   468 => (x"c8",x"86",x"70",x"98"),
   469 => (x"05",x"c6",x"87",x"c1"),
   470 => (x"cc",x"fa",x"48",x"c0"),
   471 => (x"78",x"c8",x"1e",x"c0"),
   472 => (x"e9",x"fe",x"1e",x"c1"),
   473 => (x"c5",x"d8",x"49",x"fd"),
   474 => (x"e1",x"87",x"c8",x"86"),
   475 => (x"70",x"98",x"05",x"c6"),
   476 => (x"87",x"c1",x"cc",x"fa"),
   477 => (x"48",x"c0",x"78",x"c8"),
   478 => (x"1e",x"c0",x"ea",x"c7"),
   479 => (x"1e",x"c1",x"c5",x"d8"),
   480 => (x"49",x"fd",x"c7",x"87"),
   481 => (x"c8",x"86",x"70",x"98"),
   482 => (x"05",x"c5",x"87",x"c0"),
   483 => (x"48",x"c9",x"d1",x"87"),
   484 => (x"c1",x"cc",x"fa",x"bf"),
   485 => (x"1e",x"c0",x"ea",x"d0"),
   486 => (x"1e",x"c0",x"e3",x"e3"),
   487 => (x"87",x"c8",x"86",x"c1"),
   488 => (x"cc",x"fa",x"bf",x"02"),
   489 => (x"c1",x"ed",x"87",x"c1"),
   490 => (x"c4",x"c6",x"4a",x"48"),
   491 => (x"c6",x"fe",x"a0",x"4c"),
   492 => (x"c1",x"cb",x"cc",x"bf"),
   493 => (x"4b",x"c1",x"cc",x"c4"),
   494 => (x"9f",x"bf",x"49",x"c4"),
   495 => (x"a6",x"5a",x"c5",x"d6"),
   496 => (x"ea",x"a9",x"05",x"c0"),
   497 => (x"cc",x"87",x"c8",x"a4"),
   498 => (x"4a",x"6a",x"49",x"fa"),
   499 => (x"eb",x"87",x"70",x"4b"),
   500 => (x"db",x"87",x"c7",x"fe"),
   501 => (x"a2",x"49",x"9f",x"69"),
   502 => (x"49",x"ca",x"e9",x"d5"),
   503 => (x"a9",x"02",x"c0",x"cc"),
   504 => (x"87",x"c0",x"e7",x"e5"),
   505 => (x"49",x"d6",x"fd",x"87"),
   506 => (x"c0",x"48",x"c7",x"f4"),
   507 => (x"87",x"73",x"1e",x"c0"),
   508 => (x"e8",x"c3",x"1e",x"c0"),
   509 => (x"e2",x"c9",x"87",x"c1"),
   510 => (x"c4",x"c6",x"1e",x"73"),
   511 => (x"49",x"f7",x"fa",x"87"),
   512 => (x"cc",x"86",x"70",x"98"),
   513 => (x"05",x"c0",x"c5",x"87"),
   514 => (x"c0",x"48",x"c7",x"d4"),
   515 => (x"87",x"c0",x"e8",x"db"),
   516 => (x"49",x"d6",x"d1",x"87"),
   517 => (x"c0",x"ea",x"e3",x"1e"),
   518 => (x"c0",x"e1",x"e4",x"87"),
   519 => (x"c8",x"1e",x"c0",x"ea"),
   520 => (x"fb",x"1e",x"c1",x"c5"),
   521 => (x"d8",x"49",x"fa",x"e2"),
   522 => (x"87",x"cc",x"86",x"70"),
   523 => (x"98",x"05",x"c0",x"c9"),
   524 => (x"87",x"c1",x"cc",x"ce"),
   525 => (x"48",x"c1",x"78",x"c0"),
   526 => (x"e4",x"87",x"c8",x"1e"),
   527 => (x"c0",x"eb",x"c4",x"1e"),
   528 => (x"c1",x"c4",x"fc",x"49"),
   529 => (x"fa",x"c4",x"87",x"c8"),
   530 => (x"86",x"70",x"98",x"02"),
   531 => (x"c0",x"cf",x"87",x"c0"),
   532 => (x"e9",x"c2",x"1e",x"c0"),
   533 => (x"e0",x"e9",x"87",x"c4"),
   534 => (x"86",x"c0",x"48",x"c6"),
   535 => (x"c3",x"87",x"c1",x"cc"),
   536 => (x"c4",x"97",x"bf",x"49"),
   537 => (x"c1",x"d5",x"a9",x"05"),
   538 => (x"c0",x"cd",x"87",x"c1"),
   539 => (x"cc",x"c5",x"97",x"bf"),
   540 => (x"49",x"c2",x"ea",x"a9"),
   541 => (x"02",x"c0",x"c5",x"87"),
   542 => (x"c0",x"48",x"c5",x"e4"),
   543 => (x"87",x"c1",x"c4",x"c6"),
   544 => (x"97",x"bf",x"49",x"c3"),
   545 => (x"e9",x"a9",x"02",x"c0"),
   546 => (x"d2",x"87",x"c1",x"c4"),
   547 => (x"c6",x"97",x"bf",x"49"),
   548 => (x"c3",x"eb",x"a9",x"02"),
   549 => (x"c0",x"c5",x"87",x"c0"),
   550 => (x"48",x"c5",x"c5",x"87"),
   551 => (x"c1",x"c4",x"d1",x"97"),
   552 => (x"bf",x"49",x"99",x"05"),
   553 => (x"c0",x"cc",x"87",x"c1"),
   554 => (x"c4",x"d2",x"97",x"bf"),
   555 => (x"49",x"c2",x"a9",x"02"),
   556 => (x"c0",x"c5",x"87",x"c0"),
   557 => (x"48",x"c4",x"e9",x"87"),
   558 => (x"c1",x"c4",x"d3",x"97"),
   559 => (x"bf",x"48",x"c1",x"cc"),
   560 => (x"ca",x"58",x"c1",x"88"),
   561 => (x"c1",x"cc",x"ce",x"58"),
   562 => (x"c1",x"c4",x"d4",x"97"),
   563 => (x"bf",x"49",x"73",x"81"),
   564 => (x"c1",x"c4",x"d5",x"97"),
   565 => (x"bf",x"4a",x"c8",x"32"),
   566 => (x"c1",x"cc",x"da",x"48"),
   567 => (x"72",x"a1",x"78",x"c1"),
   568 => (x"c4",x"d6",x"97",x"bf"),
   569 => (x"48",x"c1",x"cc",x"f2"),
   570 => (x"58",x"c1",x"cc",x"ce"),
   571 => (x"bf",x"02",x"c2",x"e0"),
   572 => (x"87",x"c8",x"1e",x"c0"),
   573 => (x"e9",x"df",x"1e",x"c1"),
   574 => (x"c5",x"d8",x"49",x"f7"),
   575 => (x"cd",x"87",x"c8",x"86"),
   576 => (x"70",x"98",x"02",x"c0"),
   577 => (x"c5",x"87",x"c0",x"48"),
   578 => (x"c3",x"d6",x"87",x"c1"),
   579 => (x"cc",x"c6",x"bf",x"48"),
   580 => (x"c4",x"30",x"c1",x"cc"),
   581 => (x"f6",x"58",x"c1",x"cc"),
   582 => (x"c6",x"bf",x"4a",x"c1"),
   583 => (x"cc",x"ee",x"5a",x"c1"),
   584 => (x"c4",x"eb",x"97",x"bf"),
   585 => (x"49",x"c8",x"31",x"c1"),
   586 => (x"c4",x"ea",x"97",x"bf"),
   587 => (x"4b",x"a1",x"49",x"c1"),
   588 => (x"c4",x"ec",x"97",x"bf"),
   589 => (x"4b",x"d0",x"33",x"73"),
   590 => (x"a1",x"49",x"c1",x"c4"),
   591 => (x"ed",x"97",x"bf",x"4b"),
   592 => (x"d8",x"33",x"73",x"a1"),
   593 => (x"49",x"c1",x"cc",x"fa"),
   594 => (x"59",x"c1",x"cc",x"ee"),
   595 => (x"bf",x"91",x"c1",x"cc"),
   596 => (x"da",x"bf",x"81",x"c1"),
   597 => (x"cc",x"e2",x"59",x"c1"),
   598 => (x"c4",x"f3",x"97",x"bf"),
   599 => (x"4b",x"c8",x"33",x"c1"),
   600 => (x"c4",x"f2",x"97",x"bf"),
   601 => (x"4c",x"a3",x"4b",x"c1"),
   602 => (x"c4",x"f4",x"97",x"bf"),
   603 => (x"4c",x"d0",x"34",x"74"),
   604 => (x"a3",x"4b",x"c1",x"c4"),
   605 => (x"f5",x"97",x"bf",x"4c"),
   606 => (x"cf",x"9c",x"d8",x"34"),
   607 => (x"74",x"a3",x"4b",x"c1"),
   608 => (x"cc",x"e6",x"5b",x"c2"),
   609 => (x"8b",x"73",x"92",x"c1"),
   610 => (x"cc",x"e6",x"48",x"72"),
   611 => (x"a1",x"78",x"c1",x"ce"),
   612 => (x"87",x"c1",x"c4",x"d8"),
   613 => (x"97",x"bf",x"49",x"c8"),
   614 => (x"31",x"c1",x"c4",x"d7"),
   615 => (x"97",x"bf",x"4a",x"a1"),
   616 => (x"49",x"c1",x"cc",x"f6"),
   617 => (x"59",x"c5",x"31",x"c7"),
   618 => (x"ff",x"81",x"c9",x"29"),
   619 => (x"c1",x"cc",x"ee",x"59"),
   620 => (x"c1",x"c4",x"dd",x"97"),
   621 => (x"bf",x"4a",x"c8",x"32"),
   622 => (x"c1",x"c4",x"dc",x"97"),
   623 => (x"bf",x"4b",x"a2",x"4a"),
   624 => (x"c1",x"cc",x"fa",x"5a"),
   625 => (x"c1",x"cc",x"ee",x"bf"),
   626 => (x"92",x"c1",x"cc",x"da"),
   627 => (x"bf",x"82",x"c1",x"cc"),
   628 => (x"ea",x"5a",x"c1",x"cc"),
   629 => (x"e2",x"48",x"c0",x"78"),
   630 => (x"c1",x"cc",x"de",x"48"),
   631 => (x"72",x"a1",x"78",x"c1"),
   632 => (x"48",x"26",x"f4",x"e2"),
   633 => (x"87",x"4e",x"6f",x"20"),
   634 => (x"70",x"61",x"72",x"74"),
   635 => (x"69",x"74",x"69",x"6f"),
   636 => (x"6e",x"20",x"73",x"69"),
   637 => (x"67",x"6e",x"61",x"74"),
   638 => (x"75",x"72",x"65",x"20"),
   639 => (x"66",x"6f",x"75",x"6e"),
   640 => (x"64",x"0a",x"00",x"52"),
   641 => (x"65",x"61",x"64",x"69"),
   642 => (x"6e",x"67",x"20",x"62"),
   643 => (x"6f",x"6f",x"74",x"20"),
   644 => (x"73",x"65",x"63",x"74"),
   645 => (x"6f",x"72",x"20",x"25"),
   646 => (x"64",x"0a",x"00",x"52"),
   647 => (x"65",x"61",x"64",x"20"),
   648 => (x"62",x"6f",x"6f",x"74"),
   649 => (x"20",x"73",x"65",x"63"),
   650 => (x"74",x"6f",x"72",x"20"),
   651 => (x"66",x"72",x"6f",x"6d"),
   652 => (x"20",x"66",x"69",x"72"),
   653 => (x"73",x"74",x"20",x"70"),
   654 => (x"61",x"72",x"74",x"69"),
   655 => (x"74",x"69",x"6f",x"6e"),
   656 => (x"0a",x"00",x"55",x"6e"),
   657 => (x"73",x"75",x"70",x"70"),
   658 => (x"6f",x"72",x"74",x"65"),
   659 => (x"64",x"20",x"70",x"61"),
   660 => (x"72",x"74",x"69",x"74"),
   661 => (x"69",x"6f",x"6e",x"20"),
   662 => (x"74",x"79",x"70",x"65"),
   663 => (x"21",x"0d",x"00",x"46"),
   664 => (x"41",x"54",x"33",x"32"),
   665 => (x"20",x"20",x"20",x"00"),
   666 => (x"52",x"65",x"61",x"64"),
   667 => (x"69",x"6e",x"67",x"20"),
   668 => (x"4d",x"42",x"52",x"0a"),
   669 => (x"00",x"46",x"41",x"54"),
   670 => (x"31",x"36",x"20",x"20"),
   671 => (x"20",x"00",x"46",x"41"),
   672 => (x"54",x"33",x"32",x"20"),
   673 => (x"20",x"20",x"00",x"46"),
   674 => (x"41",x"54",x"31",x"32"),
   675 => (x"20",x"20",x"20",x"00"),
   676 => (x"50",x"61",x"72",x"74"),
   677 => (x"69",x"74",x"69",x"6f"),
   678 => (x"6e",x"63",x"6f",x"75"),
   679 => (x"6e",x"74",x"20",x"25"),
   680 => (x"64",x"0a",x"00",x"48"),
   681 => (x"75",x"6e",x"74",x"69"),
   682 => (x"6e",x"67",x"20",x"66"),
   683 => (x"6f",x"72",x"20",x"66"),
   684 => (x"69",x"6c",x"65",x"73"),
   685 => (x"79",x"73",x"74",x"65"),
   686 => (x"6d",x"0a",x"00",x"46"),
   687 => (x"41",x"54",x"33",x"32"),
   688 => (x"20",x"20",x"20",x"00"),
   689 => (x"46",x"41",x"54",x"31"),
   690 => (x"36",x"20",x"20",x"20"),
   691 => (x"00",x"52",x"65",x"61"),
   692 => (x"64",x"69",x"6e",x"67"),
   693 => (x"20",x"64",x"69",x"72"),
   694 => (x"65",x"63",x"74",x"6f"),
   695 => (x"72",x"79",x"20",x"73"),
   696 => (x"65",x"63",x"74",x"6f"),
   697 => (x"72",x"20",x"25",x"64"),
   698 => (x"0a",x"00",x"66",x"69"),
   699 => (x"6c",x"65",x"20",x"22"),
   700 => (x"25",x"73",x"22",x"20"),
   701 => (x"66",x"6f",x"75",x"6e"),
   702 => (x"64",x"0d",x"00",x"47"),
   703 => (x"65",x"74",x"46",x"41"),
   704 => (x"54",x"4c",x"69",x"6e"),
   705 => (x"6b",x"20",x"72",x"65"),
   706 => (x"74",x"75",x"72",x"6e"),
   707 => (x"65",x"64",x"20",x"25"),
   708 => (x"64",x"0a",x"00",x"43"),
   709 => (x"61",x"6e",x"27",x"74"),
   710 => (x"20",x"6f",x"70",x"65"),
   711 => (x"6e",x"20",x"25",x"73"),
   712 => (x"0a",x"00",x"0e",x"5e"),
   713 => (x"5b",x"5c",x"5d",x"0e"),
   714 => (x"71",x"4a",x"c1",x"cc"),
   715 => (x"ce",x"bf",x"02",x"cc"),
   716 => (x"87",x"72",x"4b",x"c7"),
   717 => (x"b7",x"2b",x"72",x"4c"),
   718 => (x"c1",x"ff",x"9c",x"ca"),
   719 => (x"87",x"72",x"4b",x"c8"),
   720 => (x"b7",x"2b",x"72",x"4c"),
   721 => (x"c3",x"ff",x"9c",x"c1"),
   722 => (x"cc",x"fe",x"bf",x"ab"),
   723 => (x"02",x"de",x"87",x"c1"),
   724 => (x"c4",x"c6",x"1e",x"c1"),
   725 => (x"cc",x"da",x"bf",x"49"),
   726 => (x"73",x"81",x"ea",x"dd"),
   727 => (x"87",x"c4",x"86",x"70"),
   728 => (x"98",x"05",x"c5",x"87"),
   729 => (x"c0",x"48",x"c0",x"f5"),
   730 => (x"87",x"c1",x"cd",x"c2"),
   731 => (x"5b",x"c1",x"cc",x"ce"),
   732 => (x"bf",x"02",x"d8",x"87"),
   733 => (x"74",x"4a",x"c4",x"92"),
   734 => (x"c1",x"c4",x"c6",x"82"),
   735 => (x"6a",x"49",x"eb",x"f8"),
   736 => (x"87",x"70",x"49",x"4d"),
   737 => (x"cf",x"ff",x"ff",x"ff"),
   738 => (x"ff",x"9d",x"d0",x"87"),
   739 => (x"74",x"4a",x"c2",x"92"),
   740 => (x"c1",x"c4",x"c6",x"82"),
   741 => (x"9f",x"6a",x"49",x"ec"),
   742 => (x"d8",x"87",x"70",x"4d"),
   743 => (x"75",x"48",x"ed",x"e4"),
   744 => (x"87",x"0e",x"5e",x"5b"),
   745 => (x"5c",x"5d",x"0e",x"f4"),
   746 => (x"86",x"71",x"4c",x"c0"),
   747 => (x"4b",x"c1",x"cc",x"fe"),
   748 => (x"48",x"ff",x"78",x"c1"),
   749 => (x"cc",x"e2",x"bf",x"4d"),
   750 => (x"c1",x"cc",x"e6",x"bf"),
   751 => (x"7e",x"c1",x"cc",x"ce"),
   752 => (x"bf",x"02",x"c9",x"87"),
   753 => (x"c1",x"cc",x"c6",x"bf"),
   754 => (x"4a",x"c4",x"32",x"c7"),
   755 => (x"87",x"c1",x"cc",x"ea"),
   756 => (x"bf",x"4a",x"c4",x"32"),
   757 => (x"c8",x"a6",x"5a",x"c8"),
   758 => (x"a6",x"48",x"c0",x"78"),
   759 => (x"c4",x"66",x"48",x"c0"),
   760 => (x"a8",x"06",x"c3",x"cd"),
   761 => (x"87",x"c8",x"66",x"49"),
   762 => (x"cf",x"99",x"05",x"c0"),
   763 => (x"e2",x"87",x"6e",x"1e"),
   764 => (x"c0",x"eb",x"cd",x"1e"),
   765 => (x"d2",x"c9",x"87",x"c1"),
   766 => (x"c4",x"c6",x"1e",x"cc"),
   767 => (x"66",x"49",x"48",x"c1"),
   768 => (x"80",x"d0",x"a6",x"58"),
   769 => (x"71",x"e7",x"f2",x"87"),
   770 => (x"cc",x"86",x"c1",x"c4"),
   771 => (x"c6",x"4b",x"c3",x"87"),
   772 => (x"c0",x"e0",x"83",x"97"),
   773 => (x"6b",x"49",x"99",x"02"),
   774 => (x"c2",x"c5",x"87",x"97"),
   775 => (x"6b",x"49",x"c3",x"e5"),
   776 => (x"a9",x"02",x"c1",x"fb"),
   777 => (x"87",x"cb",x"a3",x"49"),
   778 => (x"97",x"69",x"49",x"d8"),
   779 => (x"99",x"05",x"c1",x"ef"),
   780 => (x"87",x"cb",x"1e",x"c0"),
   781 => (x"e0",x"66",x"1e",x"73"),
   782 => (x"49",x"ea",x"cf",x"87"),
   783 => (x"c8",x"86",x"70",x"98"),
   784 => (x"05",x"c1",x"dc",x"87"),
   785 => (x"dc",x"a3",x"4a",x"6a"),
   786 => (x"49",x"e8",x"ed",x"87"),
   787 => (x"70",x"4a",x"c4",x"a4"),
   788 => (x"49",x"72",x"79",x"da"),
   789 => (x"a3",x"4a",x"9f",x"6a"),
   790 => (x"49",x"e9",x"d6",x"87"),
   791 => (x"c4",x"a6",x"58",x"c1"),
   792 => (x"cc",x"ce",x"bf",x"02"),
   793 => (x"d8",x"87",x"d4",x"a3"),
   794 => (x"4a",x"9f",x"6a",x"49"),
   795 => (x"e9",x"c3",x"87",x"70"),
   796 => (x"49",x"c0",x"ff",x"ff"),
   797 => (x"99",x"71",x"48",x"d0"),
   798 => (x"30",x"c8",x"a6",x"58"),
   799 => (x"c5",x"87",x"c4",x"a6"),
   800 => (x"48",x"c0",x"78",x"c4"),
   801 => (x"66",x"4a",x"6e",x"82"),
   802 => (x"c8",x"a4",x"49",x"72"),
   803 => (x"79",x"c0",x"7c",x"dc"),
   804 => (x"66",x"1e",x"c0",x"eb"),
   805 => (x"ea",x"1e",x"cf",x"e7"),
   806 => (x"87",x"c8",x"86",x"c1"),
   807 => (x"48",x"c1",x"cf",x"87"),
   808 => (x"c8",x"66",x"48",x"c1"),
   809 => (x"80",x"cc",x"a6",x"58"),
   810 => (x"c8",x"66",x"48",x"c4"),
   811 => (x"66",x"a8",x"04",x"fc"),
   812 => (x"f3",x"87",x"c1",x"cc"),
   813 => (x"ce",x"bf",x"02",x"c0"),
   814 => (x"f3",x"87",x"75",x"49"),
   815 => (x"f9",x"e3",x"87",x"70"),
   816 => (x"4d",x"1e",x"c0",x"eb"),
   817 => (x"fb",x"1e",x"ce",x"f7"),
   818 => (x"87",x"c8",x"86",x"75"),
   819 => (x"49",x"cf",x"ff",x"ff"),
   820 => (x"ff",x"f8",x"99",x"a9"),
   821 => (x"02",x"d6",x"87",x"75"),
   822 => (x"49",x"c2",x"89",x"c1"),
   823 => (x"cc",x"c6",x"bf",x"91"),
   824 => (x"c1",x"cc",x"de",x"bf"),
   825 => (x"48",x"71",x"80",x"c4"),
   826 => (x"a6",x"58",x"fb",x"ea"),
   827 => (x"87",x"c0",x"48",x"f4"),
   828 => (x"8e",x"e8",x"d1",x"87"),
   829 => (x"0e",x"5e",x"5b",x"5c"),
   830 => (x"5d",x"0e",x"1e",x"71"),
   831 => (x"4b",x"1e",x"c1",x"cd"),
   832 => (x"c2",x"49",x"fa",x"dc"),
   833 => (x"87",x"c4",x"86",x"70"),
   834 => (x"98",x"02",x"c1",x"f6"),
   835 => (x"87",x"c1",x"cd",x"c6"),
   836 => (x"bf",x"49",x"c7",x"ff"),
   837 => (x"81",x"c9",x"29",x"c4"),
   838 => (x"a6",x"59",x"c0",x"4d"),
   839 => (x"4c",x"6e",x"48",x"c0"),
   840 => (x"b7",x"a8",x"06",x"c1"),
   841 => (x"ec",x"87",x"c1",x"cc"),
   842 => (x"de",x"bf",x"49",x"c1"),
   843 => (x"cd",x"ca",x"bf",x"4a"),
   844 => (x"c2",x"8a",x"c1",x"cc"),
   845 => (x"c6",x"bf",x"92",x"72"),
   846 => (x"a1",x"49",x"c1",x"cc"),
   847 => (x"ca",x"bf",x"4a",x"74"),
   848 => (x"9a",x"72",x"a1",x"49"),
   849 => (x"d4",x"66",x"1e",x"71"),
   850 => (x"e2",x"ef",x"87",x"c4"),
   851 => (x"86",x"70",x"98",x"05"),
   852 => (x"c5",x"87",x"c0",x"48"),
   853 => (x"c1",x"c0",x"87",x"c1"),
   854 => (x"84",x"c1",x"cc",x"ca"),
   855 => (x"bf",x"49",x"74",x"99"),
   856 => (x"05",x"cc",x"87",x"c1"),
   857 => (x"cd",x"ca",x"bf",x"49"),
   858 => (x"f6",x"f7",x"87",x"c1"),
   859 => (x"cd",x"ce",x"58",x"d4"),
   860 => (x"66",x"48",x"c8",x"c0"),
   861 => (x"80",x"d8",x"a6",x"58"),
   862 => (x"c1",x"85",x"6e",x"b7"),
   863 => (x"ad",x"04",x"fe",x"e5"),
   864 => (x"87",x"cf",x"87",x"73"),
   865 => (x"1e",x"c0",x"ec",x"d3"),
   866 => (x"1e",x"cb",x"f4",x"87"),
   867 => (x"c8",x"86",x"c0",x"48"),
   868 => (x"c5",x"87",x"c1",x"cd"),
   869 => (x"c6",x"bf",x"48",x"26"),
   870 => (x"e5",x"ea",x"87",x"1e"),
   871 => (x"f3",x"09",x"97",x"79"),
   872 => (x"09",x"71",x"48",x"26"),
   873 => (x"4f",x"0e",x"5e",x"5b"),
   874 => (x"5c",x"0e",x"71",x"4b"),
   875 => (x"c0",x"4c",x"13",x"4a"),
   876 => (x"9a",x"02",x"cc",x"87"),
   877 => (x"72",x"49",x"e3",x"87"),
   878 => (x"c1",x"84",x"13",x"4a"),
   879 => (x"9a",x"05",x"f4",x"87"),
   880 => (x"74",x"48",x"c2",x"87"),
   881 => (x"26",x"4d",x"26",x"4c"),
   882 => (x"26",x"4b",x"26",x"4f"),
   883 => (x"0e",x"5e",x"5b",x"5c"),
   884 => (x"5d",x"0e",x"fc",x"86"),
   885 => (x"71",x"4a",x"c0",x"e0"),
   886 => (x"66",x"4c",x"c1",x"cd"),
   887 => (x"ce",x"4b",x"c0",x"7e"),
   888 => (x"72",x"9a",x"05",x"ce"),
   889 => (x"87",x"c1",x"cd",x"cf"),
   890 => (x"4b",x"c1",x"cd",x"ce"),
   891 => (x"48",x"c0",x"f0",x"50"),
   892 => (x"c1",x"d2",x"87",x"72"),
   893 => (x"9a",x"02",x"c0",x"e9"),
   894 => (x"87",x"d4",x"66",x"4d"),
   895 => (x"72",x"1e",x"72",x"49"),
   896 => (x"75",x"4a",x"ca",x"cf"),
   897 => (x"87",x"26",x"4a",x"c0"),
   898 => (x"f9",x"f6",x"81",x"11"),
   899 => (x"53",x"71",x"1e",x"72"),
   900 => (x"49",x"75",x"4a",x"c9"),
   901 => (x"fe",x"87",x"70",x"4a"),
   902 => (x"26",x"49",x"c1",x"8c"),
   903 => (x"72",x"9a",x"05",x"ff"),
   904 => (x"da",x"87",x"c0",x"b7"),
   905 => (x"ac",x"06",x"dd",x"87"),
   906 => (x"c0",x"e4",x"66",x"02"),
   907 => (x"c5",x"87",x"c0",x"f0"),
   908 => (x"4a",x"c3",x"87",x"c0"),
   909 => (x"e0",x"4a",x"73",x"0a"),
   910 => (x"97",x"7a",x"0a",x"c1"),
   911 => (x"83",x"8c",x"c0",x"b7"),
   912 => (x"ac",x"01",x"ff",x"e3"),
   913 => (x"87",x"c1",x"cd",x"ce"),
   914 => (x"ab",x"02",x"de",x"87"),
   915 => (x"d8",x"66",x"4c",x"dc"),
   916 => (x"66",x"1e",x"c1",x"8b"),
   917 => (x"97",x"6b",x"49",x"74"),
   918 => (x"0f",x"c4",x"86",x"6e"),
   919 => (x"48",x"c1",x"80",x"c4"),
   920 => (x"a6",x"58",x"c1",x"cd"),
   921 => (x"ce",x"ab",x"05",x"ff"),
   922 => (x"e5",x"87",x"6e",x"48"),
   923 => (x"fc",x"8e",x"26",x"4d"),
   924 => (x"26",x"4c",x"26",x"4b"),
   925 => (x"26",x"4f",x"30",x"31"),
   926 => (x"32",x"33",x"34",x"35"),
   927 => (x"36",x"37",x"38",x"39"),
   928 => (x"41",x"42",x"43",x"44"),
   929 => (x"45",x"46",x"00",x"0e"),
   930 => (x"5e",x"5b",x"5c",x"5d"),
   931 => (x"0e",x"71",x"4b",x"ff"),
   932 => (x"4d",x"13",x"4c",x"74"),
   933 => (x"9c",x"02",x"d8",x"87"),
   934 => (x"c1",x"85",x"d4",x"66"),
   935 => (x"1e",x"74",x"49",x"d4"),
   936 => (x"66",x"0f",x"c4",x"86"),
   937 => (x"74",x"a8",x"05",x"c7"),
   938 => (x"87",x"13",x"4c",x"74"),
   939 => (x"9c",x"05",x"e8",x"87"),
   940 => (x"75",x"48",x"26",x"4d"),
   941 => (x"26",x"4c",x"26",x"4b"),
   942 => (x"26",x"4f",x"0e",x"5e"),
   943 => (x"5b",x"5c",x"5d",x"0e"),
   944 => (x"e8",x"86",x"c4",x"a6"),
   945 => (x"59",x"c0",x"e8",x"66"),
   946 => (x"4d",x"c0",x"4c",x"c8"),
   947 => (x"a6",x"48",x"c0",x"78"),
   948 => (x"6e",x"97",x"bf",x"4b"),
   949 => (x"6e",x"48",x"c1",x"80"),
   950 => (x"c4",x"a6",x"58",x"73"),
   951 => (x"9b",x"02",x"c6",x"d3"),
   952 => (x"87",x"c8",x"66",x"02"),
   953 => (x"c5",x"db",x"87",x"cc"),
   954 => (x"a6",x"48",x"c0",x"78"),
   955 => (x"fc",x"80",x"c0",x"78"),
   956 => (x"73",x"4a",x"c0",x"e0"),
   957 => (x"8a",x"02",x"c3",x"c6"),
   958 => (x"87",x"c3",x"8a",x"02"),
   959 => (x"c3",x"c0",x"87",x"c2"),
   960 => (x"8a",x"02",x"c2",x"e8"),
   961 => (x"87",x"c2",x"8a",x"02"),
   962 => (x"c2",x"f4",x"87",x"c4"),
   963 => (x"8a",x"02",x"c2",x"ee"),
   964 => (x"87",x"c2",x"8a",x"02"),
   965 => (x"c2",x"e8",x"87",x"c3"),
   966 => (x"8a",x"02",x"c2",x"ea"),
   967 => (x"87",x"d4",x"8a",x"02"),
   968 => (x"c0",x"f6",x"87",x"d4"),
   969 => (x"8a",x"02",x"c1",x"c0"),
   970 => (x"87",x"ca",x"8a",x"02"),
   971 => (x"c0",x"f2",x"87",x"c1"),
   972 => (x"8a",x"02",x"c1",x"e1"),
   973 => (x"87",x"c1",x"8a",x"02"),
   974 => (x"df",x"87",x"c8",x"8a"),
   975 => (x"02",x"c1",x"ce",x"87"),
   976 => (x"c4",x"8a",x"02",x"c0"),
   977 => (x"e3",x"87",x"c3",x"8a"),
   978 => (x"02",x"c0",x"e5",x"87"),
   979 => (x"c2",x"8a",x"02",x"c8"),
   980 => (x"87",x"c3",x"8a",x"02"),
   981 => (x"d3",x"87",x"c1",x"fa"),
   982 => (x"87",x"cc",x"a6",x"48"),
   983 => (x"ca",x"78",x"c2",x"d2"),
   984 => (x"87",x"cc",x"a6",x"48"),
   985 => (x"c2",x"78",x"c2",x"ca"),
   986 => (x"87",x"cc",x"a6",x"48"),
   987 => (x"d0",x"78",x"c2",x"c2"),
   988 => (x"87",x"c0",x"f0",x"66"),
   989 => (x"1e",x"c0",x"f0",x"66"),
   990 => (x"1e",x"c4",x"85",x"75"),
   991 => (x"4a",x"c4",x"8a",x"6a"),
   992 => (x"49",x"fc",x"c3",x"87"),
   993 => (x"c8",x"86",x"70",x"49"),
   994 => (x"71",x"a4",x"4c",x"c1"),
   995 => (x"e5",x"87",x"c8",x"a6"),
   996 => (x"48",x"c1",x"78",x"c1"),
   997 => (x"dd",x"87",x"c0",x"f0"),
   998 => (x"66",x"1e",x"c4",x"85"),
   999 => (x"75",x"4a",x"c4",x"8a"),
  1000 => (x"6a",x"49",x"c0",x"f0"),
  1001 => (x"66",x"0f",x"c4",x"86"),
  1002 => (x"c1",x"84",x"c1",x"c6"),
  1003 => (x"87",x"c0",x"f0",x"66"),
  1004 => (x"1e",x"c0",x"e5",x"49"),
  1005 => (x"c0",x"f0",x"66",x"0f"),
  1006 => (x"c4",x"86",x"c1",x"84"),
  1007 => (x"c0",x"f4",x"87",x"c8"),
  1008 => (x"a6",x"48",x"c1",x"78"),
  1009 => (x"c0",x"ec",x"87",x"d0"),
  1010 => (x"a6",x"48",x"c1",x"78"),
  1011 => (x"f8",x"80",x"c1",x"78"),
  1012 => (x"c0",x"e0",x"87",x"c0"),
  1013 => (x"f0",x"ab",x"06",x"da"),
  1014 => (x"87",x"c0",x"f9",x"ab"),
  1015 => (x"03",x"d4",x"87",x"d4"),
  1016 => (x"66",x"49",x"ca",x"91"),
  1017 => (x"73",x"4a",x"c0",x"f0"),
  1018 => (x"8a",x"d4",x"a6",x"48"),
  1019 => (x"72",x"a1",x"78",x"f4"),
  1020 => (x"80",x"c1",x"78",x"cc"),
  1021 => (x"66",x"02",x"c1",x"ea"),
  1022 => (x"87",x"c4",x"85",x"75"),
  1023 => (x"49",x"c4",x"89",x"a6"),
  1024 => (x"48",x"69",x"78",x"c1"),
  1025 => (x"e4",x"ab",x"05",x"d8"),
  1026 => (x"87",x"c4",x"66",x"48"),
  1027 => (x"c0",x"b7",x"a8",x"03"),
  1028 => (x"cf",x"87",x"c0",x"ed"),
  1029 => (x"49",x"f6",x"c3",x"87"),
  1030 => (x"c4",x"66",x"48",x"c0"),
  1031 => (x"08",x"88",x"c8",x"a6"),
  1032 => (x"58",x"d0",x"66",x"1e"),
  1033 => (x"d8",x"66",x"1e",x"c0"),
  1034 => (x"f8",x"66",x"1e",x"c0"),
  1035 => (x"f8",x"66",x"1e",x"dc"),
  1036 => (x"66",x"1e",x"d8",x"66"),
  1037 => (x"49",x"f6",x"d4",x"87"),
  1038 => (x"d4",x"86",x"70",x"49"),
  1039 => (x"71",x"a4",x"4c",x"c0"),
  1040 => (x"e1",x"87",x"c0",x"e5"),
  1041 => (x"ab",x"05",x"cf",x"87"),
  1042 => (x"d0",x"a6",x"48",x"c0"),
  1043 => (x"78",x"c4",x"80",x"c0"),
  1044 => (x"78",x"f4",x"80",x"c1"),
  1045 => (x"78",x"cc",x"87",x"c0"),
  1046 => (x"f0",x"66",x"1e",x"73"),
  1047 => (x"49",x"c0",x"f0",x"66"),
  1048 => (x"0f",x"c4",x"86",x"6e"),
  1049 => (x"97",x"bf",x"4b",x"6e"),
  1050 => (x"48",x"c1",x"80",x"c4"),
  1051 => (x"a6",x"58",x"73",x"9b"),
  1052 => (x"05",x"f9",x"ed",x"87"),
  1053 => (x"74",x"48",x"e8",x"8e"),
  1054 => (x"26",x"4d",x"26",x"4c"),
  1055 => (x"26",x"4b",x"26",x"4f"),
  1056 => (x"1e",x"c0",x"1e",x"c0"),
  1057 => (x"f6",x"db",x"1e",x"d0"),
  1058 => (x"a6",x"1e",x"d0",x"66"),
  1059 => (x"49",x"f8",x"ea",x"87"),
  1060 => (x"f4",x"8e",x"26",x"4f"),
  1061 => (x"1e",x"73",x"1e",x"72"),
  1062 => (x"9a",x"02",x"c0",x"e7"),
  1063 => (x"87",x"c0",x"48",x"c1"),
  1064 => (x"4b",x"72",x"a9",x"06"),
  1065 => (x"d1",x"87",x"72",x"82"),
  1066 => (x"06",x"c9",x"87",x"73"),
  1067 => (x"83",x"72",x"a9",x"01"),
  1068 => (x"f4",x"87",x"c3",x"87"),
  1069 => (x"c1",x"b2",x"3a",x"72"),
  1070 => (x"a9",x"03",x"89",x"73"),
  1071 => (x"80",x"07",x"c1",x"2a"),
  1072 => (x"2b",x"05",x"f3",x"87"),
  1073 => (x"26",x"4b",x"26",x"4f"),
  1074 => (x"1e",x"75",x"1e",x"c4"),
  1075 => (x"4d",x"71",x"b7",x"a1"),
  1076 => (x"04",x"ff",x"b9",x"c1"),
  1077 => (x"81",x"c3",x"bd",x"07"),
  1078 => (x"72",x"b7",x"a2",x"04"),
  1079 => (x"ff",x"ba",x"c1",x"82"),
  1080 => (x"c1",x"bd",x"07",x"fe"),
  1081 => (x"ee",x"87",x"c1",x"2d"),
  1082 => (x"04",x"ff",x"b8",x"c1"),
  1083 => (x"80",x"07",x"2d",x"04"),
  1084 => (x"ff",x"b9",x"c1",x"81"),
  1085 => (x"07",x"26",x"4d",x"26"),
  1086 => (x"4f",x"26",x"4d",x"26"),
	others => (others => x"00")
);

-- Xilinx XST attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "no_rw_check";

-- Altera Quartus attributes
attribute ramstyle: string;
attribute ramstyle of ram: signal is "no_rw_check";

signal q_local : word_t;
signal q2_local : word_t;

begin
    
	process(clk,q_local)
	begin

		q(31 downto 24)<=q_local(0);
		q(23 downto 16)<=q_local(1);
		q(15 downto 8)<=q_local(2);
		q(7 downto 0)<=q_local(3);

		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel(3) = '1') then
					ram(to_integer(unsigned(addr)))(3) <= d(7 downto 0);
				end if;
				if bytesel(2) = '1' then
					ram(to_integer(unsigned(addr)))(2) <= d(15 downto 8);
				end if;
				if bytesel(1) = '1' then
					ram(to_integer(unsigned(addr)))(1) <= d(23 downto 16);
				end if;
				if bytesel(0) = '1' then
					ram(to_integer(unsigned(addr)))(0) <= d(31 downto 24);
				end if;
			end if;
			q_local <= ram(to_integer(unsigned(addr)));
		end if;
	end process;

	-- Second port
	
	process(clk,q2_local)
	begin

		q2(31 downto 24)<=q2_local(0);
		q2(23 downto 16)<=q2_local(1);
		q2(15 downto 8)<=q2_local(2);
		q2(7 downto 0)<=q2_local(3);

		if(rising_edge(clk)) then 
			if(we2 = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel2(3) = '1') then
					ram(to_integer(unsigned(addr2)))(3) <= d2(7 downto 0);
				end if;
				if bytesel2(2) = '1' then
					ram(to_integer(unsigned(addr2)))(2) <= d2(15 downto 8);
				end if;
				if bytesel2(1) = '1' then
					ram(to_integer(unsigned(addr2)))(1) <= d2(23 downto 16);
				end if;
				if bytesel2(0) = '1' then
					ram(to_integer(unsigned(addr2)))(0) <= d2(31 downto 24);
				end if;
			end if;
			q2_local <= ram(to_integer(unsigned(addr2)));
		end if;
	end process;

end arch;

