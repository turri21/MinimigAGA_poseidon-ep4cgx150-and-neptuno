library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM-2 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
type ram_type is array (0 to 2 ** (maxAddrBitBRAM-3) - 1) of word_t;

signal ram : ram_type :=
(
     0 => (x"01",x"da",x"87",x"04"),
     1 => (x"dd",x"87",x"0e",x"58"),
     2 => (x"5e",x"59",x"5a",x"0e"),
     3 => (x"27",x"00",x"00",x"00"),
     4 => (x"2c",x"0f",x"26",x"4a"),
     5 => (x"26",x"49",x"26",x"48"),
     6 => (x"ff",x"80",x"26",x"08"),
     7 => (x"4f",x"27",x"00",x"00"),
     8 => (x"00",x"2d",x"4f",x"27"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"4f",x"00",x"fd",x"87"),
    11 => (x"4f",x"c1",x"ce",x"e0"),
    12 => (x"4e",x"c9",x"c0",x"86"),
    13 => (x"c1",x"ce",x"e0",x"49"),
    14 => (x"c1",x"c4",x"fc",x"48"),
    15 => (x"89",x"d0",x"89",x"03"),
    16 => (x"c0",x"40",x"40",x"40"),
    17 => (x"40",x"f6",x"87",x"d0"),
    18 => (x"81",x"05",x"c0",x"50"),
    19 => (x"c1",x"89",x"05",x"f9"),
    20 => (x"87",x"c1",x"c4",x"fc"),
    21 => (x"4d",x"c1",x"c4",x"fc"),
    22 => (x"4c",x"74",x"ad",x"02"),
    23 => (x"c4",x"87",x"24",x"0f"),
    24 => (x"f7",x"87",x"c2",x"d9"),
    25 => (x"87",x"c1",x"c4",x"fc"),
    26 => (x"4d",x"c1",x"c4",x"fc"),
    27 => (x"4c",x"74",x"ad",x"02"),
    28 => (x"c6",x"87",x"c4",x"8c"),
    29 => (x"6c",x"0f",x"f5",x"87"),
    30 => (x"00",x"fd",x"87",x"0e"),
    31 => (x"5e",x"5b",x"5c",x"0e"),
    32 => (x"c8",x"c0",x"c0",x"c0"),
    33 => (x"4b",x"c9",x"e1",x"4c"),
    34 => (x"c9",x"f3",x"bf",x"4a"),
    35 => (x"c1",x"8a",x"02",x"cb"),
    36 => (x"87",x"74",x"49",x"c1"),
    37 => (x"84",x"11",x"53",x"c1"),
    38 => (x"8a",x"05",x"f5",x"87"),
    39 => (x"c2",x"87",x"26",x"4d"),
    40 => (x"26",x"4c",x"26",x"4b"),
    41 => (x"26",x"4f",x"1e",x"73"),
    42 => (x"1e",x"71",x"4b",x"e7"),
    43 => (x"48",x"c0",x"e0",x"50"),
    44 => (x"e3",x"48",x"c8",x"50"),
    45 => (x"e3",x"48",x"c6",x"50"),
    46 => (x"e7",x"48",x"c0",x"e1"),
    47 => (x"50",x"73",x"4a",x"c8"),
    48 => (x"b7",x"2a",x"c8",x"c0"),
    49 => (x"c0",x"c0",x"49",x"ca"),
    50 => (x"81",x"71",x"0a",x"97"),
    51 => (x"7a",x"73",x"4a",x"c3"),
    52 => (x"ff",x"9a",x"c8",x"c0"),
    53 => (x"c0",x"c0",x"49",x"cb"),
    54 => (x"81",x"71",x"0a",x"97"),
    55 => (x"7a",x"e7",x"48",x"c0"),
    56 => (x"e0",x"50",x"e3",x"48"),
    57 => (x"c8",x"50",x"e3",x"48"),
    58 => (x"c0",x"50",x"e7",x"48"),
    59 => (x"c0",x"e1",x"50",x"fe"),
    60 => (x"f0",x"87",x"1e",x"73"),
    61 => (x"1e",x"c2",x"c0",x"c0"),
    62 => (x"4b",x"73",x"0f",x"fe"),
    63 => (x"e4",x"87",x"1e",x"73"),
    64 => (x"1e",x"eb",x"48",x"c3"),
    65 => (x"ef",x"50",x"e7",x"48"),
    66 => (x"c0",x"e0",x"50",x"e3"),
    67 => (x"48",x"c8",x"50",x"e3"),
    68 => (x"48",x"c6",x"50",x"e7"),
    69 => (x"48",x"c0",x"e1",x"50"),
    70 => (x"ff",x"c2",x"48",x"c1"),
    71 => (x"9f",x"78",x"e7",x"48"),
    72 => (x"c0",x"e0",x"50",x"e3"),
    73 => (x"48",x"c4",x"50",x"e3"),
    74 => (x"48",x"c2",x"50",x"e7"),
    75 => (x"48",x"c0",x"e1",x"50"),
    76 => (x"e7",x"48",x"c0",x"e0"),
    77 => (x"50",x"e3",x"48",x"c8"),
    78 => (x"50",x"e3",x"48",x"c7"),
    79 => (x"50",x"e7",x"48",x"c0"),
    80 => (x"e1",x"50",x"fc",x"f6"),
    81 => (x"87",x"c0",x"ff",x"ff"),
    82 => (x"49",x"fd",x"da",x"87"),
    83 => (x"c0",x"fc",x"c0",x"4b"),
    84 => (x"c8",x"ed",x"49",x"c0"),
    85 => (x"f2",x"cf",x"87",x"d1"),
    86 => (x"dd",x"87",x"70",x"98"),
    87 => (x"02",x"c1",x"cb",x"87"),
    88 => (x"c0",x"ff",x"f0",x"4b"),
    89 => (x"c8",x"d6",x"49",x"c0"),
    90 => (x"f1",x"fb",x"87",x"d7"),
    91 => (x"d0",x"87",x"70",x"98"),
    92 => (x"02",x"c0",x"e7",x"87"),
    93 => (x"c3",x"f0",x"4b",x"c2"),
    94 => (x"c0",x"c0",x"1e",x"c6"),
    95 => (x"fd",x"49",x"c0",x"ee"),
    96 => (x"f1",x"87",x"c4",x"86"),
    97 => (x"70",x"98",x"02",x"c9"),
    98 => (x"87",x"c3",x"ff",x"4b"),
    99 => (x"fd",x"e3",x"87",x"c0"),
   100 => (x"e0",x"87",x"c7",x"c9"),
   101 => (x"49",x"c0",x"f1",x"cd"),
   102 => (x"87",x"d7",x"87",x"c7"),
   103 => (x"de",x"49",x"c0",x"f1"),
   104 => (x"c4",x"87",x"c7",x"fa"),
   105 => (x"49",x"c0",x"f0",x"fd"),
   106 => (x"87",x"c7",x"87",x"c9"),
   107 => (x"c3",x"49",x"c0",x"f0"),
   108 => (x"f4",x"87",x"73",x"49"),
   109 => (x"fb",x"ef",x"87",x"fe"),
   110 => (x"d2",x"87",x"fb",x"e5"),
   111 => (x"87",x"38",x"33",x"32"),
   112 => (x"4f",x"53",x"44",x"41"),
   113 => (x"42",x"42",x"49",x"4e"),
   114 => (x"00",x"43",x"61",x"6e"),
   115 => (x"27",x"74",x"20",x"6c"),
   116 => (x"6f",x"61",x"64",x"20"),
   117 => (x"66",x"69",x"72",x"6d"),
   118 => (x"77",x"61",x"72",x"65"),
   119 => (x"0a",x"00",x"55",x"6e"),
   120 => (x"61",x"62",x"6c",x"65"),
   121 => (x"20",x"74",x"6f",x"20"),
   122 => (x"6c",x"6f",x"63",x"61"),
   123 => (x"74",x"65",x"20",x"70"),
   124 => (x"61",x"72",x"74",x"69"),
   125 => (x"74",x"69",x"6f",x"6e"),
   126 => (x"0a",x"00",x"55",x"6e"),
   127 => (x"61",x"62",x"6c",x"65"),
   128 => (x"20",x"74",x"6f",x"20"),
   129 => (x"6c",x"6f",x"63",x"61"),
   130 => (x"74",x"65",x"20",x"70"),
   131 => (x"61",x"72",x"74",x"69"),
   132 => (x"74",x"69",x"6f",x"6e"),
   133 => (x"0a",x"00",x"48",x"75"),
   134 => (x"6e",x"74",x"69",x"6e"),
   135 => (x"67",x"20",x"66",x"6f"),
   136 => (x"72",x"20",x"70",x"61"),
   137 => (x"72",x"74",x"69",x"74"),
   138 => (x"69",x"6f",x"6e",x"0a"),
   139 => (x"00",x"49",x"6e",x"69"),
   140 => (x"74",x"69",x"61",x"6c"),
   141 => (x"69",x"7a",x"69",x"6e"),
   142 => (x"67",x"20",x"53",x"44"),
   143 => (x"20",x"63",x"61",x"72"),
   144 => (x"64",x"0a",x"00",x"46"),
   145 => (x"61",x"69",x"6c",x"65"),
   146 => (x"64",x"20",x"74",x"6f"),
   147 => (x"20",x"69",x"6e",x"69"),
   148 => (x"74",x"69",x"61",x"6c"),
   149 => (x"69",x"7a",x"65",x"20"),
   150 => (x"53",x"44",x"20",x"63"),
   151 => (x"61",x"72",x"64",x"0a"),
   152 => (x"00",x"00",x"00",x"00"),
   153 => (x"00",x"00",x"00",x"00"),
   154 => (x"08",x"33",x"fc",x"0f"),
   155 => (x"ff",x"00",x"df",x"f1"),
   156 => (x"80",x"60",x"f6",x"00"),
   157 => (x"00",x"00",x"12",x"1e"),
   158 => (x"e4",x"86",x"e3",x"48"),
   159 => (x"c3",x"ff",x"50",x"e3"),
   160 => (x"97",x"bf",x"48",x"c4"),
   161 => (x"a6",x"58",x"6e",x"49"),
   162 => (x"c3",x"ff",x"99",x"e3"),
   163 => (x"48",x"c3",x"ff",x"50"),
   164 => (x"c8",x"31",x"e3",x"97"),
   165 => (x"bf",x"48",x"c8",x"a6"),
   166 => (x"58",x"c4",x"66",x"48"),
   167 => (x"c3",x"ff",x"98",x"cc"),
   168 => (x"a6",x"58",x"c8",x"66"),
   169 => (x"b1",x"e3",x"48",x"c3"),
   170 => (x"ff",x"50",x"c8",x"31"),
   171 => (x"e3",x"97",x"bf",x"48"),
   172 => (x"d0",x"a6",x"58",x"cc"),
   173 => (x"66",x"48",x"c3",x"ff"),
   174 => (x"98",x"d4",x"a6",x"58"),
   175 => (x"d0",x"66",x"b1",x"e3"),
   176 => (x"48",x"c3",x"ff",x"50"),
   177 => (x"c8",x"31",x"e3",x"97"),
   178 => (x"bf",x"48",x"d8",x"a6"),
   179 => (x"58",x"d4",x"66",x"48"),
   180 => (x"c3",x"ff",x"98",x"dc"),
   181 => (x"a6",x"58",x"d8",x"66"),
   182 => (x"b1",x"71",x"48",x"e4"),
   183 => (x"8e",x"26",x"4f",x"0e"),
   184 => (x"5e",x"5b",x"5c",x"0e"),
   185 => (x"1e",x"71",x"4a",x"72"),
   186 => (x"49",x"c3",x"ff",x"99"),
   187 => (x"e3",x"09",x"97",x"79"),
   188 => (x"09",x"c1",x"c4",x"fc"),
   189 => (x"bf",x"05",x"c8",x"87"),
   190 => (x"d0",x"66",x"48",x"c9"),
   191 => (x"30",x"d4",x"a6",x"58"),
   192 => (x"d0",x"66",x"49",x"d8"),
   193 => (x"29",x"c3",x"ff",x"99"),
   194 => (x"e3",x"09",x"97",x"79"),
   195 => (x"09",x"d0",x"66",x"49"),
   196 => (x"d0",x"29",x"c3",x"ff"),
   197 => (x"99",x"e3",x"09",x"97"),
   198 => (x"79",x"09",x"d0",x"66"),
   199 => (x"49",x"c8",x"29",x"c3"),
   200 => (x"ff",x"99",x"e3",x"09"),
   201 => (x"97",x"79",x"09",x"d0"),
   202 => (x"66",x"49",x"c3",x"ff"),
   203 => (x"99",x"e3",x"09",x"97"),
   204 => (x"79",x"09",x"72",x"49"),
   205 => (x"d0",x"29",x"c3",x"ff"),
   206 => (x"99",x"e3",x"09",x"97"),
   207 => (x"79",x"09",x"97",x"bf"),
   208 => (x"48",x"c4",x"a6",x"58"),
   209 => (x"6e",x"4b",x"c3",x"ff"),
   210 => (x"9b",x"c9",x"f0",x"ff"),
   211 => (x"4c",x"c3",x"ff",x"ab"),
   212 => (x"05",x"dc",x"87",x"e3"),
   213 => (x"48",x"c3",x"ff",x"50"),
   214 => (x"e3",x"97",x"bf",x"48"),
   215 => (x"c4",x"a6",x"58",x"6e"),
   216 => (x"4b",x"c3",x"ff",x"9b"),
   217 => (x"c1",x"8c",x"02",x"c6"),
   218 => (x"87",x"c3",x"ff",x"ab"),
   219 => (x"02",x"e4",x"87",x"73"),
   220 => (x"4a",x"c4",x"b7",x"2a"),
   221 => (x"c0",x"f0",x"a2",x"49"),
   222 => (x"c0",x"e9",x"e0",x"87"),
   223 => (x"73",x"4a",x"cf",x"9a"),
   224 => (x"c0",x"f0",x"a2",x"49"),
   225 => (x"c0",x"e9",x"d4",x"87"),
   226 => (x"73",x"48",x"26",x"c2"),
   227 => (x"87",x"26",x"4d",x"26"),
   228 => (x"4c",x"26",x"4b",x"26"),
   229 => (x"4f",x"1e",x"c0",x"49"),
   230 => (x"e3",x"48",x"c3",x"ff"),
   231 => (x"50",x"c1",x"81",x"c3"),
   232 => (x"c8",x"b7",x"a9",x"04"),
   233 => (x"f2",x"87",x"26",x"4f"),
   234 => (x"1e",x"73",x"1e",x"e8"),
   235 => (x"87",x"c4",x"f8",x"df"),
   236 => (x"4b",x"c0",x"1e",x"c0"),
   237 => (x"ff",x"f0",x"c1",x"f7"),
   238 => (x"49",x"fc",x"e3",x"87"),
   239 => (x"c4",x"86",x"c1",x"a8"),
   240 => (x"05",x"c0",x"e8",x"87"),
   241 => (x"e3",x"48",x"c3",x"ff"),
   242 => (x"50",x"c1",x"c0",x"c0"),
   243 => (x"c0",x"c0",x"c0",x"1e"),
   244 => (x"c0",x"e1",x"f0",x"c1"),
   245 => (x"e9",x"49",x"fc",x"c6"),
   246 => (x"87",x"c4",x"86",x"70"),
   247 => (x"98",x"05",x"c9",x"87"),
   248 => (x"e3",x"48",x"c3",x"ff"),
   249 => (x"50",x"c1",x"48",x"cb"),
   250 => (x"87",x"fe",x"e9",x"87"),
   251 => (x"c1",x"8b",x"05",x"fe"),
   252 => (x"ff",x"87",x"c0",x"48"),
   253 => (x"fe",x"da",x"87",x"43"),
   254 => (x"4d",x"44",x"34",x"31"),
   255 => (x"20",x"25",x"64",x"0a"),
   256 => (x"00",x"43",x"4d",x"44"),
   257 => (x"35",x"35",x"20",x"25"),
   258 => (x"64",x"0a",x"00",x"43"),
   259 => (x"4d",x"44",x"34",x"31"),
   260 => (x"20",x"25",x"64",x"0a"),
   261 => (x"00",x"43",x"4d",x"44"),
   262 => (x"35",x"35",x"20",x"25"),
   263 => (x"64",x"0a",x"00",x"69"),
   264 => (x"6e",x"69",x"74",x"20"),
   265 => (x"25",x"64",x"0a",x"20"),
   266 => (x"20",x"00",x"69",x"6e"),
   267 => (x"69",x"74",x"20",x"25"),
   268 => (x"64",x"0a",x"20",x"20"),
   269 => (x"00",x"43",x"6d",x"64"),
   270 => (x"5f",x"69",x"6e",x"69"),
   271 => (x"74",x"0a",x"00",x"43"),
   272 => (x"4d",x"44",x"38",x"5f"),
   273 => (x"34",x"20",x"72",x"65"),
   274 => (x"73",x"70",x"6f",x"6e"),
   275 => (x"73",x"65",x"3a",x"20"),
   276 => (x"25",x"64",x"0a",x"00"),
   277 => (x"43",x"4d",x"44",x"35"),
   278 => (x"38",x"20",x"25",x"64"),
   279 => (x"0a",x"20",x"20",x"00"),
   280 => (x"43",x"4d",x"44",x"35"),
   281 => (x"38",x"5f",x"32",x"20"),
   282 => (x"25",x"64",x"0a",x"20"),
   283 => (x"20",x"00",x"43",x"4d"),
   284 => (x"44",x"35",x"38",x"20"),
   285 => (x"25",x"64",x"0a",x"20"),
   286 => (x"20",x"00",x"53",x"44"),
   287 => (x"48",x"43",x"20",x"49"),
   288 => (x"6e",x"69",x"74",x"69"),
   289 => (x"61",x"6c",x"69",x"7a"),
   290 => (x"61",x"74",x"69",x"6f"),
   291 => (x"6e",x"20",x"65",x"72"),
   292 => (x"72",x"6f",x"72",x"21"),
   293 => (x"0a",x"00",x"63",x"6d"),
   294 => (x"64",x"5f",x"43",x"4d"),
   295 => (x"44",x"38",x"20",x"72"),
   296 => (x"65",x"73",x"70",x"6f"),
   297 => (x"6e",x"73",x"65",x"3a"),
   298 => (x"20",x"25",x"64",x"0a"),
   299 => (x"00",x"52",x"65",x"61"),
   300 => (x"64",x"20",x"63",x"6f"),
   301 => (x"6d",x"6d",x"61",x"6e"),
   302 => (x"64",x"20",x"66",x"61"),
   303 => (x"69",x"6c",x"65",x"64"),
   304 => (x"20",x"61",x"74",x"20"),
   305 => (x"25",x"64",x"20",x"28"),
   306 => (x"25",x"64",x"29",x"0a"),
   307 => (x"00",x"1e",x"73",x"1e"),
   308 => (x"e3",x"48",x"c3",x"ff"),
   309 => (x"50",x"d0",x"f5",x"49"),
   310 => (x"c0",x"e4",x"ca",x"87"),
   311 => (x"d3",x"4b",x"c0",x"1e"),
   312 => (x"c0",x"ff",x"f0",x"c1"),
   313 => (x"c1",x"49",x"f7",x"f6"),
   314 => (x"87",x"c4",x"86",x"70"),
   315 => (x"98",x"05",x"c9",x"87"),
   316 => (x"e3",x"48",x"c3",x"ff"),
   317 => (x"50",x"c1",x"48",x"cb"),
   318 => (x"87",x"fa",x"d9",x"87"),
   319 => (x"c1",x"8b",x"05",x"ff"),
   320 => (x"dc",x"87",x"c0",x"48"),
   321 => (x"fa",x"ca",x"87",x"1e"),
   322 => (x"73",x"1e",x"1e",x"fa"),
   323 => (x"c7",x"87",x"c6",x"ea"),
   324 => (x"1e",x"c0",x"e1",x"f0"),
   325 => (x"c1",x"c8",x"49",x"f7"),
   326 => (x"c5",x"87",x"70",x"4b"),
   327 => (x"73",x"1e",x"d2",x"d6"),
   328 => (x"49",x"c0",x"ee",x"de"),
   329 => (x"87",x"c8",x"86",x"c1"),
   330 => (x"ab",x"02",x"c8",x"87"),
   331 => (x"fe",x"de",x"87",x"c0"),
   332 => (x"48",x"c1",x"ff",x"87"),
   333 => (x"f5",x"c0",x"87",x"70"),
   334 => (x"49",x"cf",x"ff",x"ff"),
   335 => (x"99",x"c6",x"ea",x"a9"),
   336 => (x"02",x"c8",x"87",x"fe"),
   337 => (x"c7",x"87",x"c0",x"48"),
   338 => (x"c1",x"e8",x"87",x"e3"),
   339 => (x"48",x"c3",x"ff",x"50"),
   340 => (x"c0",x"f1",x"4b",x"f9"),
   341 => (x"d2",x"87",x"70",x"98"),
   342 => (x"02",x"c1",x"c6",x"87"),
   343 => (x"c0",x"1e",x"c0",x"ff"),
   344 => (x"f0",x"c1",x"fa",x"49"),
   345 => (x"f5",x"f8",x"87",x"c4"),
   346 => (x"86",x"70",x"98",x"05"),
   347 => (x"c0",x"f3",x"87",x"e3"),
   348 => (x"48",x"c3",x"ff",x"50"),
   349 => (x"e3",x"97",x"bf",x"48"),
   350 => (x"c4",x"a6",x"58",x"6e"),
   351 => (x"49",x"c3",x"ff",x"99"),
   352 => (x"e3",x"48",x"c3",x"ff"),
   353 => (x"50",x"e3",x"48",x"c3"),
   354 => (x"ff",x"50",x"e3",x"48"),
   355 => (x"c3",x"ff",x"50",x"e3"),
   356 => (x"48",x"c3",x"ff",x"50"),
   357 => (x"c1",x"c0",x"99",x"02"),
   358 => (x"c4",x"87",x"c1",x"48"),
   359 => (x"d5",x"87",x"c0",x"48"),
   360 => (x"d1",x"87",x"c2",x"ab"),
   361 => (x"05",x"c4",x"87",x"c0"),
   362 => (x"48",x"c8",x"87",x"c1"),
   363 => (x"8b",x"05",x"fe",x"e2"),
   364 => (x"87",x"c0",x"48",x"26"),
   365 => (x"f7",x"da",x"87",x"1e"),
   366 => (x"73",x"1e",x"c1",x"c4"),
   367 => (x"fc",x"48",x"c1",x"78"),
   368 => (x"eb",x"48",x"c3",x"ef"),
   369 => (x"50",x"c7",x"4b",x"e7"),
   370 => (x"48",x"c3",x"50",x"f7"),
   371 => (x"c7",x"87",x"e7",x"48"),
   372 => (x"c2",x"50",x"e3",x"48"),
   373 => (x"c3",x"ff",x"50",x"c0"),
   374 => (x"1e",x"c0",x"e5",x"d0"),
   375 => (x"c1",x"c0",x"49",x"f3"),
   376 => (x"fd",x"87",x"c4",x"86"),
   377 => (x"c1",x"a8",x"05",x"c2"),
   378 => (x"87",x"c1",x"4b",x"c2"),
   379 => (x"ab",x"05",x"c5",x"87"),
   380 => (x"c0",x"48",x"c0",x"f1"),
   381 => (x"87",x"c1",x"8b",x"05"),
   382 => (x"ff",x"cc",x"87",x"fc"),
   383 => (x"c9",x"87",x"c1",x"c5"),
   384 => (x"c0",x"58",x"c1",x"c4"),
   385 => (x"fc",x"bf",x"05",x"cd"),
   386 => (x"87",x"c1",x"1e",x"c0"),
   387 => (x"ff",x"f0",x"c1",x"d0"),
   388 => (x"49",x"f3",x"cb",x"87"),
   389 => (x"c4",x"86",x"e3",x"48"),
   390 => (x"c3",x"ff",x"50",x"e7"),
   391 => (x"48",x"c3",x"50",x"e3"),
   392 => (x"48",x"c3",x"ff",x"50"),
   393 => (x"c1",x"48",x"f5",x"e8"),
   394 => (x"87",x"0e",x"5e",x"5b"),
   395 => (x"5c",x"5d",x"0e",x"1e"),
   396 => (x"71",x"4a",x"c0",x"4d"),
   397 => (x"e3",x"48",x"c3",x"ff"),
   398 => (x"50",x"e7",x"48",x"c2"),
   399 => (x"50",x"eb",x"48",x"c7"),
   400 => (x"50",x"e3",x"48",x"c3"),
   401 => (x"ff",x"50",x"72",x"1e"),
   402 => (x"c0",x"ff",x"f0",x"c1"),
   403 => (x"d1",x"49",x"f2",x"ce"),
   404 => (x"87",x"c4",x"86",x"70"),
   405 => (x"98",x"05",x"c1",x"c9"),
   406 => (x"87",x"c5",x"ee",x"cd"),
   407 => (x"df",x"4b",x"e3",x"48"),
   408 => (x"c3",x"ff",x"50",x"e3"),
   409 => (x"97",x"bf",x"48",x"c4"),
   410 => (x"a6",x"58",x"6e",x"49"),
   411 => (x"c3",x"ff",x"99",x"c3"),
   412 => (x"fe",x"a9",x"05",x"de"),
   413 => (x"87",x"c0",x"4c",x"ef"),
   414 => (x"fd",x"87",x"d4",x"66"),
   415 => (x"08",x"78",x"08",x"d4"),
   416 => (x"66",x"48",x"c4",x"80"),
   417 => (x"d8",x"a6",x"58",x"c1"),
   418 => (x"84",x"c2",x"c0",x"b7"),
   419 => (x"ac",x"04",x"e7",x"87"),
   420 => (x"c1",x"4b",x"4d",x"c1"),
   421 => (x"8b",x"05",x"ff",x"c5"),
   422 => (x"87",x"e3",x"48",x"c3"),
   423 => (x"ff",x"50",x"e7",x"48"),
   424 => (x"c3",x"50",x"75",x"48"),
   425 => (x"26",x"f3",x"e5",x"87"),
   426 => (x"1e",x"73",x"1e",x"71"),
   427 => (x"4b",x"73",x"49",x"d8"),
   428 => (x"29",x"c3",x"ff",x"99"),
   429 => (x"73",x"4a",x"c8",x"2a"),
   430 => (x"cf",x"fc",x"c0",x"9a"),
   431 => (x"72",x"b1",x"73",x"4a"),
   432 => (x"c8",x"32",x"c0",x"ff"),
   433 => (x"f0",x"c0",x"c0",x"9a"),
   434 => (x"72",x"b1",x"73",x"4a"),
   435 => (x"d8",x"32",x"ff",x"c0"),
   436 => (x"c0",x"c0",x"c0",x"9a"),
   437 => (x"72",x"b1",x"71",x"48"),
   438 => (x"c4",x"87",x"26",x"4d"),
   439 => (x"26",x"4c",x"26",x"4b"),
   440 => (x"26",x"4f",x"1e",x"73"),
   441 => (x"1e",x"71",x"4b",x"73"),
   442 => (x"49",x"c8",x"29",x"c3"),
   443 => (x"ff",x"99",x"73",x"4a"),
   444 => (x"c8",x"32",x"cf",x"fc"),
   445 => (x"c0",x"9a",x"72",x"b1"),
   446 => (x"71",x"48",x"e2",x"87"),
   447 => (x"0e",x"5e",x"5b",x"5c"),
   448 => (x"0e",x"71",x"4b",x"c0"),
   449 => (x"4c",x"d0",x"66",x"48"),
   450 => (x"c0",x"b7",x"a8",x"06"),
   451 => (x"c0",x"e3",x"87",x"13"),
   452 => (x"4a",x"cc",x"66",x"97"),
   453 => (x"bf",x"49",x"cc",x"66"),
   454 => (x"48",x"c1",x"80",x"d0"),
   455 => (x"a6",x"58",x"71",x"b7"),
   456 => (x"aa",x"02",x"c4",x"87"),
   457 => (x"c1",x"48",x"cc",x"87"),
   458 => (x"c1",x"84",x"d0",x"66"),
   459 => (x"b7",x"ac",x"04",x"ff"),
   460 => (x"dd",x"87",x"c0",x"48"),
   461 => (x"c2",x"87",x"26",x"4d"),
   462 => (x"26",x"4c",x"26",x"4b"),
   463 => (x"26",x"4f",x"0e",x"5e"),
   464 => (x"5b",x"5c",x"0e",x"1e"),
   465 => (x"c1",x"cd",x"fe",x"48"),
   466 => (x"ff",x"78",x"c1",x"cd"),
   467 => (x"ce",x"48",x"c0",x"78"),
   468 => (x"c0",x"ea",x"e3",x"49"),
   469 => (x"da",x"cf",x"87",x"c1"),
   470 => (x"c5",x"c6",x"1e",x"c0"),
   471 => (x"49",x"fb",x"c9",x"87"),
   472 => (x"c4",x"86",x"70",x"98"),
   473 => (x"05",x"c5",x"87",x"c0"),
   474 => (x"48",x"ca",x"f0",x"87"),
   475 => (x"c0",x"4b",x"c1",x"cd"),
   476 => (x"fa",x"48",x"c1",x"78"),
   477 => (x"c8",x"1e",x"c0",x"ea"),
   478 => (x"f0",x"1e",x"c1",x"c5"),
   479 => (x"fc",x"49",x"fd",x"fb"),
   480 => (x"87",x"c8",x"86",x"70"),
   481 => (x"98",x"05",x"c6",x"87"),
   482 => (x"c1",x"cd",x"fa",x"48"),
   483 => (x"c0",x"78",x"c8",x"1e"),
   484 => (x"c0",x"ea",x"f9",x"1e"),
   485 => (x"c1",x"c6",x"d8",x"49"),
   486 => (x"fd",x"e1",x"87",x"c8"),
   487 => (x"86",x"70",x"98",x"05"),
   488 => (x"c6",x"87",x"c1",x"cd"),
   489 => (x"fa",x"48",x"c0",x"78"),
   490 => (x"c8",x"1e",x"c0",x"eb"),
   491 => (x"c2",x"1e",x"c1",x"c6"),
   492 => (x"d8",x"49",x"fd",x"c7"),
   493 => (x"87",x"c8",x"86",x"70"),
   494 => (x"98",x"05",x"c5",x"87"),
   495 => (x"c0",x"48",x"c9",x"db"),
   496 => (x"87",x"c1",x"cd",x"fa"),
   497 => (x"bf",x"1e",x"c0",x"eb"),
   498 => (x"cb",x"1e",x"c0",x"e3"),
   499 => (x"f5",x"87",x"c8",x"86"),
   500 => (x"c1",x"cd",x"fa",x"bf"),
   501 => (x"02",x"c1",x"ed",x"87"),
   502 => (x"c1",x"c5",x"c6",x"4a"),
   503 => (x"48",x"c6",x"fe",x"a0"),
   504 => (x"4c",x"c1",x"cc",x"cc"),
   505 => (x"bf",x"4b",x"c1",x"cd"),
   506 => (x"c4",x"9f",x"bf",x"49"),
   507 => (x"c4",x"a6",x"5a",x"c5"),
   508 => (x"d6",x"ea",x"a9",x"05"),
   509 => (x"c0",x"cc",x"87",x"c8"),
   510 => (x"a4",x"4a",x"6a",x"49"),
   511 => (x"fa",x"e9",x"87",x"70"),
   512 => (x"4b",x"db",x"87",x"c7"),
   513 => (x"fe",x"a2",x"49",x"9f"),
   514 => (x"69",x"49",x"ca",x"e9"),
   515 => (x"d5",x"a9",x"02",x"c0"),
   516 => (x"cc",x"87",x"c0",x"e8"),
   517 => (x"e0",x"49",x"d7",x"cd"),
   518 => (x"87",x"c0",x"48",x"c7"),
   519 => (x"fe",x"87",x"73",x"1e"),
   520 => (x"c0",x"e8",x"fe",x"1e"),
   521 => (x"c0",x"e2",x"db",x"87"),
   522 => (x"c1",x"c5",x"c6",x"1e"),
   523 => (x"73",x"49",x"f7",x"f8"),
   524 => (x"87",x"cc",x"86",x"70"),
   525 => (x"98",x"05",x"c0",x"c5"),
   526 => (x"87",x"c0",x"48",x"c7"),
   527 => (x"de",x"87",x"c0",x"e9"),
   528 => (x"d6",x"49",x"d6",x"e1"),
   529 => (x"87",x"c0",x"eb",x"de"),
   530 => (x"1e",x"c0",x"e1",x"f6"),
   531 => (x"87",x"c8",x"1e",x"c0"),
   532 => (x"eb",x"f6",x"1e",x"c1"),
   533 => (x"c6",x"d8",x"49",x"fa"),
   534 => (x"e2",x"87",x"cc",x"86"),
   535 => (x"70",x"98",x"05",x"c0"),
   536 => (x"c9",x"87",x"c1",x"cd"),
   537 => (x"ce",x"48",x"c1",x"78"),
   538 => (x"c0",x"e4",x"87",x"c8"),
   539 => (x"1e",x"c0",x"eb",x"ff"),
   540 => (x"1e",x"c1",x"c5",x"fc"),
   541 => (x"49",x"fa",x"c4",x"87"),
   542 => (x"c8",x"86",x"70",x"98"),
   543 => (x"02",x"c0",x"cf",x"87"),
   544 => (x"c0",x"e9",x"fd",x"1e"),
   545 => (x"c0",x"e0",x"fb",x"87"),
   546 => (x"c4",x"86",x"c0",x"48"),
   547 => (x"c6",x"cd",x"87",x"c1"),
   548 => (x"cd",x"c4",x"97",x"bf"),
   549 => (x"49",x"c1",x"d5",x"a9"),
   550 => (x"05",x"c0",x"cd",x"87"),
   551 => (x"c1",x"cd",x"c5",x"97"),
   552 => (x"bf",x"49",x"c2",x"ea"),
   553 => (x"a9",x"02",x"c0",x"c5"),
   554 => (x"87",x"c0",x"48",x"c5"),
   555 => (x"ee",x"87",x"c1",x"c5"),
   556 => (x"c6",x"97",x"bf",x"49"),
   557 => (x"c3",x"e9",x"a9",x"02"),
   558 => (x"c0",x"d2",x"87",x"c1"),
   559 => (x"c5",x"c6",x"97",x"bf"),
   560 => (x"49",x"c3",x"eb",x"a9"),
   561 => (x"02",x"c0",x"c5",x"87"),
   562 => (x"c0",x"48",x"c5",x"cf"),
   563 => (x"87",x"c1",x"c5",x"d1"),
   564 => (x"97",x"bf",x"49",x"71"),
   565 => (x"99",x"05",x"c0",x"cc"),
   566 => (x"87",x"c1",x"c5",x"d2"),
   567 => (x"97",x"bf",x"49",x"c2"),
   568 => (x"a9",x"02",x"c0",x"c5"),
   569 => (x"87",x"c0",x"48",x"c4"),
   570 => (x"f2",x"87",x"c1",x"c5"),
   571 => (x"d3",x"97",x"bf",x"48"),
   572 => (x"c1",x"cd",x"ca",x"58"),
   573 => (x"c1",x"cd",x"c6",x"bf"),
   574 => (x"48",x"c1",x"88",x"c1"),
   575 => (x"cd",x"ce",x"58",x"c1"),
   576 => (x"c5",x"d4",x"97",x"bf"),
   577 => (x"49",x"73",x"81",x"c1"),
   578 => (x"c5",x"d5",x"97",x"bf"),
   579 => (x"4a",x"c8",x"32",x"c1"),
   580 => (x"cd",x"da",x"48",x"72"),
   581 => (x"a1",x"78",x"c1",x"c5"),
   582 => (x"d6",x"97",x"bf",x"48"),
   583 => (x"c1",x"cd",x"f2",x"58"),
   584 => (x"c1",x"cd",x"ce",x"bf"),
   585 => (x"02",x"c2",x"e2",x"87"),
   586 => (x"c8",x"1e",x"c0",x"ea"),
   587 => (x"da",x"1e",x"c1",x"c6"),
   588 => (x"d8",x"49",x"f7",x"c7"),
   589 => (x"87",x"c8",x"86",x"70"),
   590 => (x"98",x"02",x"c0",x"c5"),
   591 => (x"87",x"c0",x"48",x"c3"),
   592 => (x"da",x"87",x"c1",x"cd"),
   593 => (x"c6",x"bf",x"48",x"c4"),
   594 => (x"30",x"c1",x"cd",x"f6"),
   595 => (x"58",x"c1",x"cd",x"c6"),
   596 => (x"bf",x"4a",x"c1",x"cd"),
   597 => (x"ee",x"5a",x"c1",x"c5"),
   598 => (x"eb",x"97",x"bf",x"49"),
   599 => (x"c8",x"31",x"c1",x"c5"),
   600 => (x"ea",x"97",x"bf",x"4b"),
   601 => (x"73",x"a1",x"49",x"c1"),
   602 => (x"c5",x"ec",x"97",x"bf"),
   603 => (x"4b",x"d0",x"33",x"73"),
   604 => (x"a1",x"49",x"c1",x"c5"),
   605 => (x"ed",x"97",x"bf",x"4b"),
   606 => (x"d8",x"33",x"73",x"a1"),
   607 => (x"49",x"c1",x"cd",x"fa"),
   608 => (x"59",x"c1",x"cd",x"ee"),
   609 => (x"bf",x"91",x"c1",x"cd"),
   610 => (x"da",x"bf",x"81",x"c1"),
   611 => (x"cd",x"e2",x"59",x"c1"),
   612 => (x"c5",x"f3",x"97",x"bf"),
   613 => (x"4b",x"c8",x"33",x"c1"),
   614 => (x"c5",x"f2",x"97",x"bf"),
   615 => (x"4c",x"74",x"a3",x"4b"),
   616 => (x"c1",x"c5",x"f4",x"97"),
   617 => (x"bf",x"4c",x"d0",x"34"),
   618 => (x"74",x"a3",x"4b",x"c1"),
   619 => (x"c5",x"f5",x"97",x"bf"),
   620 => (x"4c",x"cf",x"9c",x"d8"),
   621 => (x"34",x"74",x"a3",x"4b"),
   622 => (x"c1",x"cd",x"e6",x"5b"),
   623 => (x"c2",x"8b",x"73",x"92"),
   624 => (x"c1",x"cd",x"e6",x"48"),
   625 => (x"72",x"a1",x"78",x"c1"),
   626 => (x"d0",x"87",x"c1",x"c5"),
   627 => (x"d8",x"97",x"bf",x"49"),
   628 => (x"c8",x"31",x"c1",x"c5"),
   629 => (x"d7",x"97",x"bf",x"4a"),
   630 => (x"72",x"a1",x"49",x"c1"),
   631 => (x"cd",x"f6",x"59",x"c5"),
   632 => (x"31",x"c7",x"ff",x"81"),
   633 => (x"c9",x"29",x"c1",x"cd"),
   634 => (x"ee",x"59",x"c1",x"c5"),
   635 => (x"dd",x"97",x"bf",x"4a"),
   636 => (x"c8",x"32",x"c1",x"c5"),
   637 => (x"dc",x"97",x"bf",x"4b"),
   638 => (x"73",x"a2",x"4a",x"c1"),
   639 => (x"cd",x"fa",x"5a",x"c1"),
   640 => (x"cd",x"ee",x"bf",x"92"),
   641 => (x"c1",x"cd",x"da",x"bf"),
   642 => (x"82",x"c1",x"cd",x"ea"),
   643 => (x"5a",x"c1",x"cd",x"e2"),
   644 => (x"48",x"c0",x"78",x"c1"),
   645 => (x"cd",x"de",x"48",x"72"),
   646 => (x"a1",x"78",x"c1",x"48"),
   647 => (x"26",x"f4",x"d8",x"87"),
   648 => (x"4e",x"6f",x"20",x"70"),
   649 => (x"61",x"72",x"74",x"69"),
   650 => (x"74",x"69",x"6f",x"6e"),
   651 => (x"20",x"73",x"69",x"67"),
   652 => (x"6e",x"61",x"74",x"75"),
   653 => (x"72",x"65",x"20",x"66"),
   654 => (x"6f",x"75",x"6e",x"64"),
   655 => (x"0a",x"00",x"52",x"65"),
   656 => (x"61",x"64",x"69",x"6e"),
   657 => (x"67",x"20",x"62",x"6f"),
   658 => (x"6f",x"74",x"20",x"73"),
   659 => (x"65",x"63",x"74",x"6f"),
   660 => (x"72",x"20",x"25",x"64"),
   661 => (x"0a",x"00",x"52",x"65"),
   662 => (x"61",x"64",x"20",x"62"),
   663 => (x"6f",x"6f",x"74",x"20"),
   664 => (x"73",x"65",x"63",x"74"),
   665 => (x"6f",x"72",x"20",x"66"),
   666 => (x"72",x"6f",x"6d",x"20"),
   667 => (x"66",x"69",x"72",x"73"),
   668 => (x"74",x"20",x"70",x"61"),
   669 => (x"72",x"74",x"69",x"74"),
   670 => (x"69",x"6f",x"6e",x"0a"),
   671 => (x"00",x"55",x"6e",x"73"),
   672 => (x"75",x"70",x"70",x"6f"),
   673 => (x"72",x"74",x"65",x"64"),
   674 => (x"20",x"70",x"61",x"72"),
   675 => (x"74",x"69",x"74",x"69"),
   676 => (x"6f",x"6e",x"20",x"74"),
   677 => (x"79",x"70",x"65",x"21"),
   678 => (x"0d",x"00",x"46",x"41"),
   679 => (x"54",x"33",x"32",x"20"),
   680 => (x"20",x"20",x"00",x"52"),
   681 => (x"65",x"61",x"64",x"69"),
   682 => (x"6e",x"67",x"20",x"4d"),
   683 => (x"42",x"52",x"0a",x"00"),
   684 => (x"46",x"41",x"54",x"31"),
   685 => (x"36",x"20",x"20",x"20"),
   686 => (x"00",x"46",x"41",x"54"),
   687 => (x"33",x"32",x"20",x"20"),
   688 => (x"20",x"00",x"46",x"41"),
   689 => (x"54",x"31",x"32",x"20"),
   690 => (x"20",x"20",x"00",x"50"),
   691 => (x"61",x"72",x"74",x"69"),
   692 => (x"74",x"69",x"6f",x"6e"),
   693 => (x"63",x"6f",x"75",x"6e"),
   694 => (x"74",x"20",x"25",x"64"),
   695 => (x"0a",x"00",x"48",x"75"),
   696 => (x"6e",x"74",x"69",x"6e"),
   697 => (x"67",x"20",x"66",x"6f"),
   698 => (x"72",x"20",x"66",x"69"),
   699 => (x"6c",x"65",x"73",x"79"),
   700 => (x"73",x"74",x"65",x"6d"),
   701 => (x"0a",x"00",x"46",x"41"),
   702 => (x"54",x"33",x"32",x"20"),
   703 => (x"20",x"20",x"00",x"46"),
   704 => (x"41",x"54",x"31",x"36"),
   705 => (x"20",x"20",x"20",x"00"),
   706 => (x"52",x"65",x"61",x"64"),
   707 => (x"69",x"6e",x"67",x"20"),
   708 => (x"64",x"69",x"72",x"65"),
   709 => (x"63",x"74",x"6f",x"72"),
   710 => (x"79",x"20",x"73",x"65"),
   711 => (x"63",x"74",x"6f",x"72"),
   712 => (x"20",x"25",x"64",x"0a"),
   713 => (x"00",x"66",x"69",x"6c"),
   714 => (x"65",x"20",x"22",x"25"),
   715 => (x"73",x"22",x"20",x"66"),
   716 => (x"6f",x"75",x"6e",x"64"),
   717 => (x"0d",x"00",x"47",x"65"),
   718 => (x"74",x"46",x"41",x"54"),
   719 => (x"4c",x"69",x"6e",x"6b"),
   720 => (x"20",x"72",x"65",x"74"),
   721 => (x"75",x"72",x"6e",x"65"),
   722 => (x"64",x"20",x"25",x"64"),
   723 => (x"0a",x"00",x"43",x"61"),
   724 => (x"6e",x"27",x"74",x"20"),
   725 => (x"6f",x"70",x"65",x"6e"),
   726 => (x"20",x"25",x"73",x"0a"),
   727 => (x"00",x"0e",x"5e",x"5b"),
   728 => (x"5c",x"5d",x"0e",x"71"),
   729 => (x"4a",x"c1",x"cd",x"ce"),
   730 => (x"bf",x"02",x"cc",x"87"),
   731 => (x"72",x"4b",x"c7",x"b7"),
   732 => (x"2b",x"72",x"4c",x"c1"),
   733 => (x"ff",x"9c",x"ca",x"87"),
   734 => (x"72",x"4b",x"c8",x"b7"),
   735 => (x"2b",x"72",x"4c",x"c3"),
   736 => (x"ff",x"9c",x"c1",x"cd"),
   737 => (x"fe",x"bf",x"ab",x"02"),
   738 => (x"de",x"87",x"c1",x"c5"),
   739 => (x"c6",x"1e",x"c1",x"cd"),
   740 => (x"da",x"bf",x"49",x"73"),
   741 => (x"81",x"ea",x"d1",x"87"),
   742 => (x"c4",x"86",x"70",x"98"),
   743 => (x"05",x"c5",x"87",x"c0"),
   744 => (x"48",x"c0",x"f6",x"87"),
   745 => (x"c1",x"ce",x"c2",x"5b"),
   746 => (x"c1",x"cd",x"ce",x"bf"),
   747 => (x"02",x"d9",x"87",x"74"),
   748 => (x"4a",x"c4",x"92",x"c1"),
   749 => (x"c5",x"c6",x"82",x"6a"),
   750 => (x"49",x"eb",x"ec",x"87"),
   751 => (x"70",x"49",x"71",x"4d"),
   752 => (x"cf",x"ff",x"ff",x"ff"),
   753 => (x"ff",x"9d",x"d0",x"87"),
   754 => (x"74",x"4a",x"c2",x"92"),
   755 => (x"c1",x"c5",x"c6",x"82"),
   756 => (x"9f",x"6a",x"49",x"ec"),
   757 => (x"cc",x"87",x"70",x"4d"),
   758 => (x"75",x"48",x"ed",x"d9"),
   759 => (x"87",x"0e",x"5e",x"5b"),
   760 => (x"5c",x"5d",x"0e",x"f4"),
   761 => (x"86",x"71",x"4c",x"c0"),
   762 => (x"4b",x"c1",x"cd",x"fe"),
   763 => (x"48",x"ff",x"78",x"c1"),
   764 => (x"cd",x"e2",x"bf",x"4d"),
   765 => (x"c1",x"cd",x"e6",x"bf"),
   766 => (x"7e",x"c1",x"cd",x"ce"),
   767 => (x"bf",x"02",x"c9",x"87"),
   768 => (x"c1",x"cd",x"c6",x"bf"),
   769 => (x"4a",x"c4",x"32",x"c7"),
   770 => (x"87",x"c1",x"cd",x"ea"),
   771 => (x"bf",x"4a",x"c4",x"32"),
   772 => (x"c8",x"a6",x"5a",x"c8"),
   773 => (x"a6",x"48",x"c0",x"78"),
   774 => (x"c4",x"66",x"48",x"c0"),
   775 => (x"a8",x"06",x"c3",x"cf"),
   776 => (x"87",x"c8",x"66",x"49"),
   777 => (x"cf",x"99",x"05",x"c0"),
   778 => (x"e3",x"87",x"6e",x"1e"),
   779 => (x"c0",x"ec",x"c8",x"1e"),
   780 => (x"d2",x"d0",x"87",x"c1"),
   781 => (x"c5",x"c6",x"1e",x"cc"),
   782 => (x"66",x"49",x"48",x"c1"),
   783 => (x"80",x"d0",x"a6",x"58"),
   784 => (x"71",x"49",x"e7",x"e4"),
   785 => (x"87",x"cc",x"86",x"c1"),
   786 => (x"c5",x"c6",x"4b",x"c3"),
   787 => (x"87",x"c0",x"e0",x"83"),
   788 => (x"97",x"6b",x"49",x"71"),
   789 => (x"99",x"02",x"c2",x"c5"),
   790 => (x"87",x"97",x"6b",x"49"),
   791 => (x"c3",x"e5",x"a9",x"02"),
   792 => (x"c1",x"fb",x"87",x"cb"),
   793 => (x"a3",x"49",x"97",x"69"),
   794 => (x"49",x"d8",x"99",x"05"),
   795 => (x"c1",x"ef",x"87",x"cb"),
   796 => (x"1e",x"c0",x"e0",x"66"),
   797 => (x"1e",x"73",x"49",x"ea"),
   798 => (x"c2",x"87",x"c8",x"86"),
   799 => (x"70",x"98",x"05",x"c1"),
   800 => (x"dc",x"87",x"dc",x"a3"),
   801 => (x"4a",x"6a",x"49",x"e8"),
   802 => (x"de",x"87",x"70",x"4a"),
   803 => (x"c4",x"a4",x"49",x"72"),
   804 => (x"79",x"da",x"a3",x"4a"),
   805 => (x"9f",x"6a",x"49",x"e9"),
   806 => (x"c8",x"87",x"c4",x"a6"),
   807 => (x"58",x"c1",x"cd",x"ce"),
   808 => (x"bf",x"02",x"d8",x"87"),
   809 => (x"d4",x"a3",x"4a",x"9f"),
   810 => (x"6a",x"49",x"e8",x"f5"),
   811 => (x"87",x"70",x"49",x"c0"),
   812 => (x"ff",x"ff",x"99",x"71"),
   813 => (x"48",x"d0",x"30",x"c8"),
   814 => (x"a6",x"58",x"c5",x"87"),
   815 => (x"c4",x"a6",x"48",x"c0"),
   816 => (x"78",x"c4",x"66",x"4a"),
   817 => (x"6e",x"82",x"c8",x"a4"),
   818 => (x"49",x"72",x"79",x"c0"),
   819 => (x"7c",x"dc",x"66",x"1e"),
   820 => (x"c0",x"ec",x"e5",x"1e"),
   821 => (x"cf",x"ec",x"87",x"c8"),
   822 => (x"86",x"c1",x"48",x"c1"),
   823 => (x"d0",x"87",x"c8",x"66"),
   824 => (x"48",x"c1",x"80",x"cc"),
   825 => (x"a6",x"58",x"c8",x"66"),
   826 => (x"48",x"c4",x"66",x"a8"),
   827 => (x"04",x"fc",x"f1",x"87"),
   828 => (x"c1",x"cd",x"ce",x"bf"),
   829 => (x"02",x"c0",x"f4",x"87"),
   830 => (x"75",x"49",x"f9",x"e0"),
   831 => (x"87",x"70",x"4d",x"75"),
   832 => (x"1e",x"c0",x"ec",x"f6"),
   833 => (x"1e",x"ce",x"fb",x"87"),
   834 => (x"c8",x"86",x"75",x"49"),
   835 => (x"cf",x"ff",x"ff",x"ff"),
   836 => (x"f8",x"99",x"a9",x"02"),
   837 => (x"d6",x"87",x"75",x"49"),
   838 => (x"c2",x"89",x"c1",x"cd"),
   839 => (x"c6",x"bf",x"91",x"c1"),
   840 => (x"cd",x"de",x"bf",x"48"),
   841 => (x"71",x"80",x"c4",x"a6"),
   842 => (x"58",x"fb",x"e7",x"87"),
   843 => (x"c0",x"48",x"f4",x"8e"),
   844 => (x"e8",x"c3",x"87",x"0e"),
   845 => (x"5e",x"5b",x"5c",x"5d"),
   846 => (x"0e",x"1e",x"71",x"4b"),
   847 => (x"73",x"1e",x"c1",x"ce"),
   848 => (x"c2",x"49",x"fa",x"d8"),
   849 => (x"87",x"c4",x"86",x"70"),
   850 => (x"98",x"02",x"c1",x"f7"),
   851 => (x"87",x"c1",x"ce",x"c6"),
   852 => (x"bf",x"49",x"c7",x"ff"),
   853 => (x"81",x"c9",x"29",x"c4"),
   854 => (x"a6",x"59",x"c0",x"4d"),
   855 => (x"4c",x"6e",x"48",x"c0"),
   856 => (x"b7",x"a8",x"06",x"c1"),
   857 => (x"ed",x"87",x"c1",x"cd"),
   858 => (x"de",x"bf",x"49",x"c1"),
   859 => (x"ce",x"ca",x"bf",x"4a"),
   860 => (x"c2",x"8a",x"c1",x"cd"),
   861 => (x"c6",x"bf",x"92",x"72"),
   862 => (x"a1",x"49",x"c1",x"cd"),
   863 => (x"ca",x"bf",x"4a",x"74"),
   864 => (x"9a",x"72",x"a1",x"49"),
   865 => (x"d4",x"66",x"1e",x"71"),
   866 => (x"49",x"e2",x"dd",x"87"),
   867 => (x"c4",x"86",x"70",x"98"),
   868 => (x"05",x"c5",x"87",x"c0"),
   869 => (x"48",x"c1",x"c0",x"87"),
   870 => (x"c1",x"84",x"c1",x"cd"),
   871 => (x"ca",x"bf",x"49",x"74"),
   872 => (x"99",x"05",x"cc",x"87"),
   873 => (x"c1",x"ce",x"ca",x"bf"),
   874 => (x"49",x"f6",x"f1",x"87"),
   875 => (x"c1",x"ce",x"ce",x"58"),
   876 => (x"d4",x"66",x"48",x"c8"),
   877 => (x"c0",x"80",x"d8",x"a6"),
   878 => (x"58",x"c1",x"85",x"6e"),
   879 => (x"b7",x"ad",x"04",x"fe"),
   880 => (x"e4",x"87",x"cf",x"87"),
   881 => (x"73",x"1e",x"c0",x"ed"),
   882 => (x"ce",x"1e",x"cb",x"f6"),
   883 => (x"87",x"c8",x"86",x"c0"),
   884 => (x"48",x"c5",x"87",x"c1"),
   885 => (x"ce",x"c6",x"bf",x"48"),
   886 => (x"26",x"e5",x"da",x"87"),
   887 => (x"1e",x"f3",x"09",x"97"),
   888 => (x"79",x"09",x"71",x"48"),
   889 => (x"26",x"4f",x"0e",x"5e"),
   890 => (x"5b",x"5c",x"0e",x"71"),
   891 => (x"4b",x"c0",x"4c",x"13"),
   892 => (x"4a",x"72",x"9a",x"02"),
   893 => (x"cd",x"87",x"72",x"49"),
   894 => (x"e2",x"87",x"c1",x"84"),
   895 => (x"13",x"4a",x"72",x"9a"),
   896 => (x"05",x"f3",x"87",x"74"),
   897 => (x"48",x"c2",x"87",x"26"),
   898 => (x"4d",x"26",x"4c",x"26"),
   899 => (x"4b",x"26",x"4f",x"0e"),
   900 => (x"5e",x"5b",x"5c",x"5d"),
   901 => (x"0e",x"fc",x"86",x"71"),
   902 => (x"4a",x"c0",x"e0",x"66"),
   903 => (x"4c",x"c1",x"ce",x"ce"),
   904 => (x"4b",x"c0",x"7e",x"72"),
   905 => (x"9a",x"05",x"ce",x"87"),
   906 => (x"c1",x"ce",x"cf",x"4b"),
   907 => (x"c1",x"ce",x"ce",x"48"),
   908 => (x"c0",x"f0",x"50",x"c1"),
   909 => (x"d2",x"87",x"72",x"9a"),
   910 => (x"02",x"c0",x"e9",x"87"),
   911 => (x"d4",x"66",x"4d",x"72"),
   912 => (x"1e",x"72",x"49",x"75"),
   913 => (x"4a",x"ca",x"cf",x"87"),
   914 => (x"26",x"4a",x"c0",x"fa"),
   915 => (x"f9",x"81",x"11",x"53"),
   916 => (x"71",x"1e",x"72",x"49"),
   917 => (x"75",x"4a",x"c9",x"fe"),
   918 => (x"87",x"70",x"4a",x"26"),
   919 => (x"49",x"c1",x"8c",x"72"),
   920 => (x"9a",x"05",x"ff",x"da"),
   921 => (x"87",x"c0",x"b7",x"ac"),
   922 => (x"06",x"dd",x"87",x"c0"),
   923 => (x"e4",x"66",x"02",x"c5"),
   924 => (x"87",x"c0",x"f0",x"4a"),
   925 => (x"c3",x"87",x"c0",x"e0"),
   926 => (x"4a",x"73",x"0a",x"97"),
   927 => (x"7a",x"0a",x"c1",x"83"),
   928 => (x"8c",x"c0",x"b7",x"ac"),
   929 => (x"01",x"ff",x"e3",x"87"),
   930 => (x"c1",x"ce",x"ce",x"ab"),
   931 => (x"02",x"de",x"87",x"d8"),
   932 => (x"66",x"4c",x"dc",x"66"),
   933 => (x"1e",x"c1",x"8b",x"97"),
   934 => (x"6b",x"49",x"74",x"0f"),
   935 => (x"c4",x"86",x"6e",x"48"),
   936 => (x"c1",x"80",x"c4",x"a6"),
   937 => (x"58",x"c1",x"ce",x"ce"),
   938 => (x"ab",x"05",x"ff",x"e5"),
   939 => (x"87",x"6e",x"48",x"fc"),
   940 => (x"8e",x"26",x"4d",x"26"),
   941 => (x"4c",x"26",x"4b",x"26"),
   942 => (x"4f",x"30",x"31",x"32"),
   943 => (x"33",x"34",x"35",x"36"),
   944 => (x"37",x"38",x"39",x"41"),
   945 => (x"42",x"43",x"44",x"45"),
   946 => (x"46",x"00",x"0e",x"5e"),
   947 => (x"5b",x"5c",x"5d",x"0e"),
   948 => (x"71",x"4b",x"ff",x"4d"),
   949 => (x"13",x"4c",x"74",x"9c"),
   950 => (x"02",x"d8",x"87",x"c1"),
   951 => (x"85",x"d4",x"66",x"1e"),
   952 => (x"74",x"49",x"d4",x"66"),
   953 => (x"0f",x"c4",x"86",x"74"),
   954 => (x"a8",x"05",x"c7",x"87"),
   955 => (x"13",x"4c",x"74",x"9c"),
   956 => (x"05",x"e8",x"87",x"75"),
   957 => (x"48",x"26",x"4d",x"26"),
   958 => (x"4c",x"26",x"4b",x"26"),
   959 => (x"4f",x"0e",x"5e",x"5b"),
   960 => (x"5c",x"5d",x"0e",x"e8"),
   961 => (x"86",x"c4",x"a6",x"59"),
   962 => (x"c0",x"e8",x"66",x"4d"),
   963 => (x"c0",x"4c",x"c8",x"a6"),
   964 => (x"48",x"c0",x"78",x"6e"),
   965 => (x"97",x"bf",x"4b",x"6e"),
   966 => (x"48",x"c1",x"80",x"c4"),
   967 => (x"a6",x"58",x"73",x"9b"),
   968 => (x"02",x"c6",x"d3",x"87"),
   969 => (x"c8",x"66",x"02",x"c5"),
   970 => (x"db",x"87",x"cc",x"a6"),
   971 => (x"48",x"c0",x"78",x"fc"),
   972 => (x"80",x"c0",x"78",x"73"),
   973 => (x"4a",x"c0",x"e0",x"8a"),
   974 => (x"02",x"c3",x"c6",x"87"),
   975 => (x"c3",x"8a",x"02",x"c3"),
   976 => (x"c0",x"87",x"c2",x"8a"),
   977 => (x"02",x"c2",x"e8",x"87"),
   978 => (x"c2",x"8a",x"02",x"c2"),
   979 => (x"f4",x"87",x"c4",x"8a"),
   980 => (x"02",x"c2",x"ee",x"87"),
   981 => (x"c2",x"8a",x"02",x"c2"),
   982 => (x"e8",x"87",x"c3",x"8a"),
   983 => (x"02",x"c2",x"ea",x"87"),
   984 => (x"d4",x"8a",x"02",x"c0"),
   985 => (x"f6",x"87",x"d4",x"8a"),
   986 => (x"02",x"c1",x"c0",x"87"),
   987 => (x"ca",x"8a",x"02",x"c0"),
   988 => (x"f2",x"87",x"c1",x"8a"),
   989 => (x"02",x"c1",x"e1",x"87"),
   990 => (x"c1",x"8a",x"02",x"df"),
   991 => (x"87",x"c8",x"8a",x"02"),
   992 => (x"c1",x"ce",x"87",x"c4"),
   993 => (x"8a",x"02",x"c0",x"e3"),
   994 => (x"87",x"c3",x"8a",x"02"),
   995 => (x"c0",x"e5",x"87",x"c2"),
   996 => (x"8a",x"02",x"c8",x"87"),
   997 => (x"c3",x"8a",x"02",x"d3"),
   998 => (x"87",x"c1",x"fa",x"87"),
   999 => (x"cc",x"a6",x"48",x"ca"),
  1000 => (x"78",x"c2",x"d2",x"87"),
  1001 => (x"cc",x"a6",x"48",x"c2"),
  1002 => (x"78",x"c2",x"ca",x"87"),
  1003 => (x"cc",x"a6",x"48",x"d0"),
  1004 => (x"78",x"c2",x"c2",x"87"),
  1005 => (x"c0",x"f0",x"66",x"1e"),
  1006 => (x"c0",x"f0",x"66",x"1e"),
  1007 => (x"c4",x"85",x"75",x"4a"),
  1008 => (x"c4",x"8a",x"6a",x"49"),
  1009 => (x"fc",x"c3",x"87",x"c8"),
  1010 => (x"86",x"70",x"49",x"71"),
  1011 => (x"a4",x"4c",x"c1",x"e5"),
  1012 => (x"87",x"c8",x"a6",x"48"),
  1013 => (x"c1",x"78",x"c1",x"dd"),
  1014 => (x"87",x"c0",x"f0",x"66"),
  1015 => (x"1e",x"c4",x"85",x"75"),
  1016 => (x"4a",x"c4",x"8a",x"6a"),
  1017 => (x"49",x"c0",x"f0",x"66"),
  1018 => (x"0f",x"c4",x"86",x"c1"),
  1019 => (x"84",x"c1",x"c6",x"87"),
  1020 => (x"c0",x"f0",x"66",x"1e"),
  1021 => (x"c0",x"e5",x"49",x"c0"),
  1022 => (x"f0",x"66",x"0f",x"c4"),
  1023 => (x"86",x"c1",x"84",x"c0"),
  1024 => (x"f4",x"87",x"c8",x"a6"),
  1025 => (x"48",x"c1",x"78",x"c0"),
  1026 => (x"ec",x"87",x"d0",x"a6"),
  1027 => (x"48",x"c1",x"78",x"f8"),
  1028 => (x"80",x"c1",x"78",x"c0"),
  1029 => (x"e0",x"87",x"c0",x"f0"),
  1030 => (x"ab",x"06",x"da",x"87"),
  1031 => (x"c0",x"f9",x"ab",x"03"),
  1032 => (x"d4",x"87",x"d4",x"66"),
  1033 => (x"49",x"ca",x"91",x"73"),
  1034 => (x"4a",x"c0",x"f0",x"8a"),
  1035 => (x"d4",x"a6",x"48",x"72"),
  1036 => (x"a1",x"78",x"f4",x"80"),
  1037 => (x"c1",x"78",x"cc",x"66"),
  1038 => (x"02",x"c1",x"ea",x"87"),
  1039 => (x"c4",x"85",x"75",x"49"),
  1040 => (x"c4",x"89",x"a6",x"48"),
  1041 => (x"69",x"78",x"c1",x"e4"),
  1042 => (x"ab",x"05",x"d8",x"87"),
  1043 => (x"c4",x"66",x"48",x"c0"),
  1044 => (x"b7",x"a8",x"03",x"cf"),
  1045 => (x"87",x"c0",x"ed",x"49"),
  1046 => (x"f6",x"c1",x"87",x"c4"),
  1047 => (x"66",x"48",x"c0",x"08"),
  1048 => (x"88",x"c8",x"a6",x"58"),
  1049 => (x"d0",x"66",x"1e",x"d8"),
  1050 => (x"66",x"1e",x"c0",x"f8"),
  1051 => (x"66",x"1e",x"c0",x"f8"),
  1052 => (x"66",x"1e",x"dc",x"66"),
  1053 => (x"1e",x"d8",x"66",x"49"),
  1054 => (x"f6",x"d4",x"87",x"d4"),
  1055 => (x"86",x"70",x"49",x"71"),
  1056 => (x"a4",x"4c",x"c0",x"e1"),
  1057 => (x"87",x"c0",x"e5",x"ab"),
  1058 => (x"05",x"cf",x"87",x"d0"),
  1059 => (x"a6",x"48",x"c0",x"78"),
  1060 => (x"c4",x"80",x"c0",x"78"),
  1061 => (x"f4",x"80",x"c1",x"78"),
  1062 => (x"cc",x"87",x"c0",x"f0"),
  1063 => (x"66",x"1e",x"73",x"49"),
  1064 => (x"c0",x"f0",x"66",x"0f"),
  1065 => (x"c4",x"86",x"6e",x"97"),
  1066 => (x"bf",x"4b",x"6e",x"48"),
  1067 => (x"c1",x"80",x"c4",x"a6"),
  1068 => (x"58",x"73",x"9b",x"05"),
  1069 => (x"f9",x"ed",x"87",x"74"),
  1070 => (x"48",x"e8",x"8e",x"26"),
  1071 => (x"4d",x"26",x"4c",x"26"),
  1072 => (x"4b",x"26",x"4f",x"1e"),
  1073 => (x"c0",x"1e",x"c0",x"f7"),
  1074 => (x"dc",x"1e",x"d0",x"a6"),
  1075 => (x"1e",x"d0",x"66",x"49"),
  1076 => (x"f8",x"ea",x"87",x"f4"),
  1077 => (x"8e",x"26",x"4f",x"1e"),
  1078 => (x"73",x"1e",x"72",x"9a"),
  1079 => (x"02",x"c0",x"e7",x"87"),
  1080 => (x"c0",x"48",x"c1",x"4b"),
  1081 => (x"72",x"a9",x"06",x"d1"),
  1082 => (x"87",x"72",x"82",x"06"),
  1083 => (x"c9",x"87",x"73",x"83"),
  1084 => (x"72",x"a9",x"01",x"f4"),
  1085 => (x"87",x"c3",x"87",x"c1"),
  1086 => (x"b2",x"3a",x"72",x"a9"),
  1087 => (x"03",x"89",x"73",x"80"),
  1088 => (x"07",x"c1",x"2a",x"2b"),
  1089 => (x"05",x"f3",x"87",x"26"),
  1090 => (x"4b",x"26",x"4f",x"1e"),
  1091 => (x"75",x"1e",x"c4",x"4d"),
  1092 => (x"71",x"b7",x"a1",x"04"),
  1093 => (x"ff",x"b9",x"c1",x"81"),
  1094 => (x"c3",x"bd",x"07",x"72"),
  1095 => (x"b7",x"a2",x"04",x"ff"),
  1096 => (x"ba",x"c1",x"82",x"c1"),
  1097 => (x"bd",x"07",x"fe",x"ee"),
  1098 => (x"87",x"c1",x"2d",x"04"),
  1099 => (x"ff",x"b8",x"c1",x"80"),
  1100 => (x"07",x"2d",x"04",x"ff"),
  1101 => (x"b9",x"c1",x"81",x"07"),
  1102 => (x"26",x"4d",x"26",x"4f"),
	others => (others => x"00")
);

-- Xilinx XST attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "no_rw_check";

-- Altera Quartus attributes
attribute ramstyle: string;
attribute ramstyle of ram: signal is "no_rw_check";

signal q_local : word_t;

begin
    
	process(clk,q_local)
	begin

		q(31 downto 24)<=q_local(0);
		q(23 downto 16)<=q_local(1);
		q(15 downto 8)<=q_local(2);
		q(7 downto 0)<=q_local(3);

		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel(3) = '1') then
					ram(to_integer(unsigned(addr)))(3) <= d(7 downto 0);
				end if;
				if bytesel(2) = '1' then
					ram(to_integer(unsigned(addr)))(2) <= d(15 downto 8);
				end if;
				if bytesel(1) = '1' then
					ram(to_integer(unsigned(addr)))(1) <= d(23 downto 16);
				end if;
				if bytesel(0) = '1' then
					ram(to_integer(unsigned(addr)))(0) <= d(31 downto 24);
				end if;
			end if;
			q_local <= ram(to_integer(unsigned(addr)));
		end if;
	end process;

end arch;

