library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM-2 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111";
	-- Second port
	addr2 : in std_logic_vector(maxAddrBitBRAM-2 downto 0) := (others=>'0');
	q2 : out std_logic_vector(31 downto 0);
	d2 : in std_logic_vector(31 downto 0) := X"00000000";
	we2 : in std_logic := '0';
	bytesel2 : in std_logic_vector(3 downto 0) := "1111"	
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
type ram_type is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

signal ram : ram_type :=
(
     0 => (x"01",x"da",x"87",x"04"),
     1 => (x"dd",x"87",x"0e",x"58"),
     2 => (x"5e",x"59",x"5a",x"0e"),
     3 => (x"27",x"00",x"00",x"00"),
     4 => (x"29",x"0f",x"26",x"4a"),
     5 => (x"26",x"49",x"26",x"48"),
     6 => (x"ff",x"80",x"26",x"08"),
     7 => (x"4f",x"27",x"00",x"00"),
     8 => (x"00",x"2d",x"4f",x"27"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"4f",x"4f",x"00",x"fd"),
    11 => (x"87",x"c1",x"cc",x"fc"),
    12 => (x"4e",x"c9",x"c0",x"48"),
    13 => (x"c2",x"28",x"c1",x"d5"),
    14 => (x"ea",x"e5",x"d6",x"ea"),
    15 => (x"49",x"71",x"46",x"c1"),
    16 => (x"88",x"01",x"f9",x"87"),
    17 => (x"c1",x"cc",x"fc",x"49"),
    18 => (x"c1",x"c3",x"d8",x"48"),
    19 => (x"89",x"d0",x"89",x"03"),
    20 => (x"c0",x"40",x"40",x"40"),
    21 => (x"40",x"f6",x"87",x"d0"),
    22 => (x"81",x"05",x"c0",x"50"),
    23 => (x"c1",x"89",x"05",x"f9"),
    24 => (x"87",x"c1",x"c3",x"d8"),
    25 => (x"4d",x"c1",x"c3",x"d8"),
    26 => (x"4c",x"74",x"ad",x"02"),
    27 => (x"c4",x"87",x"24",x"0f"),
    28 => (x"f7",x"87",x"c2",x"db"),
    29 => (x"87",x"c1",x"c3",x"d8"),
    30 => (x"4d",x"c1",x"c3",x"d8"),
    31 => (x"4c",x"74",x"ad",x"02"),
    32 => (x"c6",x"87",x"c4",x"8c"),
    33 => (x"6c",x"0f",x"f5",x"87"),
    34 => (x"00",x"fd",x"87",x"0e"),
    35 => (x"5e",x"5b",x"5c",x"0e"),
    36 => (x"c4",x"c0",x"c0",x"c0"),
    37 => (x"4b",x"c9",x"cf",x"4c"),
    38 => (x"c9",x"e1",x"bf",x"4a"),
    39 => (x"49",x"c1",x"8a",x"71"),
    40 => (x"99",x"02",x"cf",x"87"),
    41 => (x"74",x"49",x"c1",x"84"),
    42 => (x"11",x"53",x"72",x"49"),
    43 => (x"c1",x"8a",x"71",x"99"),
    44 => (x"05",x"f1",x"87",x"c2"),
    45 => (x"87",x"26",x"4d",x"26"),
    46 => (x"4c",x"26",x"4b",x"26"),
    47 => (x"4f",x"1e",x"73",x"1e"),
    48 => (x"71",x"4b",x"e7",x"48"),
    49 => (x"c0",x"e0",x"50",x"e3"),
    50 => (x"48",x"c8",x"50",x"e3"),
    51 => (x"48",x"c6",x"50",x"e7"),
    52 => (x"48",x"c0",x"e1",x"50"),
    53 => (x"73",x"4a",x"c8",x"b7"),
    54 => (x"2a",x"c4",x"c0",x"c0"),
    55 => (x"c0",x"49",x"ca",x"81"),
    56 => (x"72",x"51",x"73",x"4a"),
    57 => (x"c3",x"ff",x"9a",x"c4"),
    58 => (x"c0",x"c0",x"c0",x"49"),
    59 => (x"cb",x"81",x"72",x"51"),
    60 => (x"e7",x"48",x"c0",x"e0"),
    61 => (x"50",x"e3",x"48",x"c8"),
    62 => (x"50",x"e3",x"48",x"c0"),
    63 => (x"50",x"e7",x"48",x"c0"),
    64 => (x"e1",x"50",x"fe",x"f4"),
    65 => (x"87",x"1e",x"73",x"1e"),
    66 => (x"c2",x"c0",x"c0",x"4b"),
    67 => (x"0f",x"fe",x"e9",x"87"),
    68 => (x"1e",x"73",x"1e",x"eb"),
    69 => (x"48",x"c3",x"ef",x"50"),
    70 => (x"e7",x"48",x"c0",x"e0"),
    71 => (x"50",x"e3",x"48",x"c8"),
    72 => (x"50",x"e3",x"48",x"c6"),
    73 => (x"50",x"e7",x"48",x"c0"),
    74 => (x"e1",x"50",x"ff",x"c2"),
    75 => (x"48",x"c1",x"9f",x"78"),
    76 => (x"e7",x"48",x"c0",x"e0"),
    77 => (x"50",x"e3",x"48",x"c4"),
    78 => (x"50",x"e3",x"48",x"c2"),
    79 => (x"50",x"e7",x"48",x"c0"),
    80 => (x"e1",x"50",x"e7",x"48"),
    81 => (x"c0",x"e0",x"50",x"e3"),
    82 => (x"48",x"c8",x"50",x"e3"),
    83 => (x"48",x"c7",x"50",x"e7"),
    84 => (x"48",x"c0",x"e1",x"50"),
    85 => (x"fc",x"f4",x"87",x"c0"),
    86 => (x"ff",x"ff",x"49",x"fd"),
    87 => (x"df",x"87",x"c0",x"fc"),
    88 => (x"c0",x"4b",x"c8",x"db"),
    89 => (x"49",x"c0",x"f0",x"ed"),
    90 => (x"87",x"d0",x"da",x"87"),
    91 => (x"70",x"98",x"02",x"c1"),
    92 => (x"c3",x"87",x"c0",x"ff"),
    93 => (x"f0",x"4b",x"c8",x"c4"),
    94 => (x"49",x"c0",x"f0",x"d9"),
    95 => (x"87",x"d6",x"c4",x"87"),
    96 => (x"70",x"98",x"02",x"c0"),
    97 => (x"e6",x"87",x"c3",x"f0"),
    98 => (x"4b",x"c2",x"c0",x"c0"),
    99 => (x"1e",x"c7",x"c7",x"49"),
   100 => (x"c0",x"ed",x"d4",x"87"),
   101 => (x"c4",x"86",x"70",x"98"),
   102 => (x"02",x"c8",x"87",x"c3"),
   103 => (x"ff",x"4b",x"fd",x"e4"),
   104 => (x"87",x"d9",x"87",x"c7"),
   105 => (x"d3",x"49",x"c0",x"ef"),
   106 => (x"ec",x"87",x"d0",x"87"),
   107 => (x"c7",x"e8",x"49",x"c0"),
   108 => (x"ef",x"e3",x"87",x"c7"),
   109 => (x"87",x"c8",x"f1",x"49"),
   110 => (x"c0",x"ef",x"da",x"87"),
   111 => (x"73",x"49",x"fb",x"fc"),
   112 => (x"87",x"fe",x"da",x"87"),
   113 => (x"fb",x"f2",x"87",x"38"),
   114 => (x"33",x"32",x"4f",x"53"),
   115 => (x"44",x"41",x"44",x"42"),
   116 => (x"49",x"4e",x"00",x"43"),
   117 => (x"61",x"6e",x"27",x"74"),
   118 => (x"20",x"6c",x"6f",x"61"),
   119 => (x"64",x"20",x"66",x"69"),
   120 => (x"72",x"6d",x"77",x"61"),
   121 => (x"72",x"65",x"0a",x"00"),
   122 => (x"55",x"6e",x"61",x"62"),
   123 => (x"6c",x"65",x"20",x"74"),
   124 => (x"6f",x"20",x"6c",x"6f"),
   125 => (x"63",x"61",x"74",x"65"),
   126 => (x"20",x"70",x"61",x"72"),
   127 => (x"74",x"69",x"74",x"69"),
   128 => (x"6f",x"6e",x"0a",x"00"),
   129 => (x"48",x"75",x"6e",x"74"),
   130 => (x"69",x"6e",x"67",x"20"),
   131 => (x"66",x"6f",x"72",x"20"),
   132 => (x"70",x"61",x"72",x"74"),
   133 => (x"69",x"74",x"69",x"6f"),
   134 => (x"6e",x"0a",x"00",x"49"),
   135 => (x"6e",x"69",x"74",x"69"),
   136 => (x"61",x"6c",x"69",x"7a"),
   137 => (x"69",x"6e",x"67",x"20"),
   138 => (x"53",x"44",x"20",x"63"),
   139 => (x"61",x"72",x"64",x"0a"),
   140 => (x"00",x"46",x"61",x"69"),
   141 => (x"6c",x"65",x"64",x"20"),
   142 => (x"74",x"6f",x"20",x"69"),
   143 => (x"6e",x"69",x"74",x"69"),
   144 => (x"61",x"6c",x"69",x"7a"),
   145 => (x"65",x"20",x"53",x"44"),
   146 => (x"20",x"63",x"61",x"72"),
   147 => (x"64",x"0a",x"00",x"00"),
   148 => (x"00",x"00",x"00",x"00"),
   149 => (x"00",x"00",x"08",x"33"),
   150 => (x"fc",x"0f",x"ff",x"00"),
   151 => (x"df",x"f1",x"80",x"60"),
   152 => (x"f6",x"00",x"00",x"00"),
   153 => (x"12",x"1e",x"e4",x"86"),
   154 => (x"e3",x"48",x"c3",x"ff"),
   155 => (x"50",x"e3",x"97",x"bf"),
   156 => (x"7e",x"6e",x"49",x"c3"),
   157 => (x"ff",x"99",x"e3",x"48"),
   158 => (x"c3",x"ff",x"50",x"c8"),
   159 => (x"31",x"e3",x"97",x"bf"),
   160 => (x"48",x"c8",x"a6",x"58"),
   161 => (x"c3",x"ff",x"98",x"cc"),
   162 => (x"a6",x"58",x"70",x"b1"),
   163 => (x"e3",x"48",x"c3",x"ff"),
   164 => (x"50",x"c8",x"31",x"e3"),
   165 => (x"97",x"bf",x"48",x"d0"),
   166 => (x"a6",x"58",x"c3",x"ff"),
   167 => (x"98",x"d4",x"a6",x"58"),
   168 => (x"70",x"b1",x"e3",x"48"),
   169 => (x"c3",x"ff",x"50",x"c8"),
   170 => (x"31",x"e3",x"97",x"bf"),
   171 => (x"48",x"d8",x"a6",x"58"),
   172 => (x"c3",x"ff",x"98",x"dc"),
   173 => (x"a6",x"58",x"70",x"b1"),
   174 => (x"71",x"48",x"e4",x"8e"),
   175 => (x"26",x"4f",x"0e",x"5e"),
   176 => (x"5b",x"5c",x"0e",x"1e"),
   177 => (x"71",x"4a",x"49",x"c3"),
   178 => (x"ff",x"99",x"e3",x"48"),
   179 => (x"71",x"50",x"c1",x"c3"),
   180 => (x"d8",x"bf",x"05",x"c8"),
   181 => (x"87",x"d0",x"66",x"48"),
   182 => (x"c9",x"30",x"d4",x"a6"),
   183 => (x"58",x"d0",x"66",x"49"),
   184 => (x"d8",x"29",x"c3",x"ff"),
   185 => (x"99",x"e3",x"48",x"71"),
   186 => (x"50",x"d0",x"66",x"49"),
   187 => (x"d0",x"29",x"c3",x"ff"),
   188 => (x"99",x"e3",x"48",x"71"),
   189 => (x"50",x"d0",x"66",x"49"),
   190 => (x"c8",x"29",x"c3",x"ff"),
   191 => (x"99",x"e3",x"48",x"71"),
   192 => (x"50",x"d0",x"66",x"49"),
   193 => (x"c3",x"ff",x"99",x"e3"),
   194 => (x"48",x"71",x"50",x"72"),
   195 => (x"49",x"d0",x"29",x"c3"),
   196 => (x"ff",x"99",x"e3",x"48"),
   197 => (x"71",x"50",x"e3",x"97"),
   198 => (x"bf",x"7e",x"6e",x"4b"),
   199 => (x"c3",x"ff",x"9b",x"c9"),
   200 => (x"f0",x"ff",x"4c",x"c3"),
   201 => (x"ff",x"ab",x"05",x"d9"),
   202 => (x"87",x"e3",x"48",x"c3"),
   203 => (x"ff",x"50",x"e3",x"97"),
   204 => (x"bf",x"7e",x"6e",x"4b"),
   205 => (x"c3",x"ff",x"9b",x"c1"),
   206 => (x"8c",x"02",x"c6",x"87"),
   207 => (x"c3",x"ff",x"ab",x"02"),
   208 => (x"e7",x"87",x"73",x"4a"),
   209 => (x"c4",x"b7",x"2a",x"c0"),
   210 => (x"f0",x"a2",x"49",x"c0"),
   211 => (x"e8",x"ff",x"87",x"73"),
   212 => (x"4a",x"cf",x"9a",x"c0"),
   213 => (x"f0",x"a2",x"49",x"c0"),
   214 => (x"e8",x"f3",x"87",x"73"),
   215 => (x"48",x"26",x"c2",x"87"),
   216 => (x"26",x"4d",x"26",x"4c"),
   217 => (x"26",x"4b",x"26",x"4f"),
   218 => (x"1e",x"c0",x"49",x"e3"),
   219 => (x"48",x"c3",x"ff",x"50"),
   220 => (x"c1",x"81",x"c3",x"c8"),
   221 => (x"b7",x"a9",x"04",x"f2"),
   222 => (x"87",x"26",x"4f",x"1e"),
   223 => (x"73",x"1e",x"e8",x"87"),
   224 => (x"c4",x"f8",x"df",x"4b"),
   225 => (x"c0",x"1e",x"c0",x"ff"),
   226 => (x"f0",x"c1",x"f7",x"49"),
   227 => (x"fc",x"ef",x"87",x"c4"),
   228 => (x"86",x"c1",x"a8",x"05"),
   229 => (x"c0",x"e8",x"87",x"e3"),
   230 => (x"48",x"c3",x"ff",x"50"),
   231 => (x"c1",x"c0",x"c0",x"c0"),
   232 => (x"c0",x"c0",x"1e",x"c0"),
   233 => (x"e1",x"f0",x"c1",x"e9"),
   234 => (x"49",x"fc",x"d2",x"87"),
   235 => (x"c4",x"86",x"70",x"98"),
   236 => (x"05",x"c9",x"87",x"e3"),
   237 => (x"48",x"c3",x"ff",x"50"),
   238 => (x"c1",x"48",x"cb",x"87"),
   239 => (x"fe",x"e9",x"87",x"c1"),
   240 => (x"8b",x"05",x"fe",x"ff"),
   241 => (x"87",x"c0",x"48",x"fe"),
   242 => (x"da",x"87",x"43",x"4d"),
   243 => (x"44",x"34",x"31",x"20"),
   244 => (x"25",x"64",x"0a",x"00"),
   245 => (x"43",x"4d",x"44",x"35"),
   246 => (x"35",x"20",x"25",x"64"),
   247 => (x"0a",x"00",x"43",x"4d"),
   248 => (x"44",x"34",x"31",x"20"),
   249 => (x"25",x"64",x"0a",x"00"),
   250 => (x"43",x"4d",x"44",x"35"),
   251 => (x"35",x"20",x"25",x"64"),
   252 => (x"0a",x"00",x"69",x"6e"),
   253 => (x"69",x"74",x"20",x"25"),
   254 => (x"64",x"0a",x"20",x"20"),
   255 => (x"00",x"69",x"6e",x"69"),
   256 => (x"74",x"20",x"25",x"64"),
   257 => (x"0a",x"20",x"20",x"00"),
   258 => (x"43",x"6d",x"64",x"5f"),
   259 => (x"69",x"6e",x"69",x"74"),
   260 => (x"0a",x"00",x"43",x"4d"),
   261 => (x"44",x"38",x"5f",x"34"),
   262 => (x"20",x"72",x"65",x"73"),
   263 => (x"70",x"6f",x"6e",x"73"),
   264 => (x"65",x"3a",x"20",x"25"),
   265 => (x"64",x"0a",x"00",x"43"),
   266 => (x"4d",x"44",x"35",x"38"),
   267 => (x"20",x"25",x"64",x"0a"),
   268 => (x"20",x"20",x"00",x"43"),
   269 => (x"4d",x"44",x"35",x"38"),
   270 => (x"5f",x"32",x"20",x"25"),
   271 => (x"64",x"0a",x"20",x"20"),
   272 => (x"00",x"43",x"4d",x"44"),
   273 => (x"35",x"38",x"20",x"25"),
   274 => (x"64",x"0a",x"20",x"20"),
   275 => (x"00",x"53",x"44",x"48"),
   276 => (x"43",x"20",x"49",x"6e"),
   277 => (x"69",x"74",x"69",x"61"),
   278 => (x"6c",x"69",x"7a",x"61"),
   279 => (x"74",x"69",x"6f",x"6e"),
   280 => (x"20",x"65",x"72",x"72"),
   281 => (x"6f",x"72",x"21",x"0a"),
   282 => (x"00",x"63",x"6d",x"64"),
   283 => (x"5f",x"43",x"4d",x"44"),
   284 => (x"38",x"20",x"72",x"65"),
   285 => (x"73",x"70",x"6f",x"6e"),
   286 => (x"73",x"65",x"3a",x"20"),
   287 => (x"25",x"64",x"0a",x"00"),
   288 => (x"52",x"65",x"61",x"64"),
   289 => (x"20",x"63",x"6f",x"6d"),
   290 => (x"6d",x"61",x"6e",x"64"),
   291 => (x"20",x"66",x"61",x"69"),
   292 => (x"6c",x"65",x"64",x"20"),
   293 => (x"61",x"74",x"20",x"25"),
   294 => (x"64",x"20",x"28",x"25"),
   295 => (x"64",x"29",x"0a",x"00"),
   296 => (x"1e",x"73",x"1e",x"e3"),
   297 => (x"48",x"c3",x"ff",x"50"),
   298 => (x"d0",x"c8",x"49",x"c0"),
   299 => (x"e3",x"e7",x"87",x"d3"),
   300 => (x"4b",x"c0",x"1e",x"c0"),
   301 => (x"ff",x"f0",x"c1",x"c1"),
   302 => (x"49",x"f8",x"c2",x"87"),
   303 => (x"c4",x"86",x"70",x"98"),
   304 => (x"05",x"c9",x"87",x"e3"),
   305 => (x"48",x"c3",x"ff",x"50"),
   306 => (x"c1",x"48",x"cb",x"87"),
   307 => (x"fa",x"d9",x"87",x"c1"),
   308 => (x"8b",x"05",x"ff",x"dc"),
   309 => (x"87",x"c0",x"48",x"fa"),
   310 => (x"ca",x"87",x"1e",x"73"),
   311 => (x"1e",x"1e",x"fa",x"c7"),
   312 => (x"87",x"c6",x"ea",x"1e"),
   313 => (x"c0",x"e1",x"f0",x"c1"),
   314 => (x"c8",x"49",x"f7",x"d1"),
   315 => (x"87",x"70",x"4b",x"1e"),
   316 => (x"d1",x"e9",x"1e",x"c0"),
   317 => (x"ed",x"e8",x"87",x"cc"),
   318 => (x"86",x"c1",x"ab",x"02"),
   319 => (x"c8",x"87",x"fe",x"df"),
   320 => (x"87",x"c0",x"48",x"c1"),
   321 => (x"fc",x"87",x"f5",x"dc"),
   322 => (x"87",x"70",x"49",x"cf"),
   323 => (x"ff",x"ff",x"99",x"c6"),
   324 => (x"ea",x"a9",x"02",x"c8"),
   325 => (x"87",x"fe",x"c8",x"87"),
   326 => (x"c0",x"48",x"c1",x"e5"),
   327 => (x"87",x"e3",x"48",x"c3"),
   328 => (x"ff",x"50",x"c0",x"f1"),
   329 => (x"4b",x"f9",x"d3",x"87"),
   330 => (x"70",x"98",x"02",x"c1"),
   331 => (x"c3",x"87",x"c0",x"1e"),
   332 => (x"c0",x"ff",x"f0",x"c1"),
   333 => (x"fa",x"49",x"f6",x"c5"),
   334 => (x"87",x"c4",x"86",x"70"),
   335 => (x"98",x"05",x"c0",x"f0"),
   336 => (x"87",x"e3",x"48",x"c3"),
   337 => (x"ff",x"50",x"e3",x"97"),
   338 => (x"bf",x"7e",x"6e",x"49"),
   339 => (x"c3",x"ff",x"99",x"e3"),
   340 => (x"48",x"c3",x"ff",x"50"),
   341 => (x"e3",x"48",x"c3",x"ff"),
   342 => (x"50",x"e3",x"48",x"c3"),
   343 => (x"ff",x"50",x"e3",x"48"),
   344 => (x"c3",x"ff",x"50",x"c1"),
   345 => (x"c0",x"99",x"02",x"c4"),
   346 => (x"87",x"c1",x"48",x"d5"),
   347 => (x"87",x"c0",x"48",x"d1"),
   348 => (x"87",x"c2",x"ab",x"05"),
   349 => (x"c4",x"87",x"c0",x"48"),
   350 => (x"c8",x"87",x"c1",x"8b"),
   351 => (x"05",x"fe",x"e5",x"87"),
   352 => (x"c0",x"48",x"26",x"f7"),
   353 => (x"de",x"87",x"1e",x"73"),
   354 => (x"1e",x"c1",x"c3",x"d8"),
   355 => (x"48",x"c1",x"78",x"eb"),
   356 => (x"48",x"c3",x"ef",x"50"),
   357 => (x"c7",x"4b",x"e7",x"48"),
   358 => (x"c3",x"50",x"f7",x"cb"),
   359 => (x"87",x"e7",x"48",x"c2"),
   360 => (x"50",x"e3",x"48",x"c3"),
   361 => (x"ff",x"50",x"c0",x"1e"),
   362 => (x"c0",x"e5",x"d0",x"c1"),
   363 => (x"c0",x"49",x"f4",x"cd"),
   364 => (x"87",x"c4",x"86",x"c1"),
   365 => (x"a8",x"05",x"c1",x"87"),
   366 => (x"4b",x"c2",x"ab",x"05"),
   367 => (x"c5",x"87",x"c0",x"48"),
   368 => (x"c0",x"ef",x"87",x"c1"),
   369 => (x"8b",x"05",x"ff",x"cd"),
   370 => (x"87",x"fc",x"ce",x"87"),
   371 => (x"c1",x"c3",x"dc",x"58"),
   372 => (x"70",x"98",x"05",x"cd"),
   373 => (x"87",x"c1",x"1e",x"c0"),
   374 => (x"ff",x"f0",x"c1",x"d0"),
   375 => (x"49",x"f3",x"de",x"87"),
   376 => (x"c4",x"86",x"e3",x"48"),
   377 => (x"c3",x"ff",x"50",x"e7"),
   378 => (x"48",x"c3",x"50",x"e3"),
   379 => (x"48",x"c3",x"ff",x"50"),
   380 => (x"c1",x"48",x"f5",x"ef"),
   381 => (x"87",x"0e",x"5e",x"5b"),
   382 => (x"5c",x"5d",x"0e",x"1e"),
   383 => (x"71",x"4a",x"c0",x"4d"),
   384 => (x"e3",x"48",x"c3",x"ff"),
   385 => (x"50",x"e7",x"48",x"c2"),
   386 => (x"50",x"eb",x"48",x"c7"),
   387 => (x"50",x"e3",x"48",x"c3"),
   388 => (x"ff",x"50",x"72",x"1e"),
   389 => (x"c0",x"ff",x"f0",x"c1"),
   390 => (x"d1",x"49",x"f2",x"e1"),
   391 => (x"87",x"c4",x"86",x"70"),
   392 => (x"98",x"05",x"c1",x"c5"),
   393 => (x"87",x"c5",x"ee",x"cd"),
   394 => (x"df",x"4b",x"e3",x"48"),
   395 => (x"c3",x"ff",x"50",x"e3"),
   396 => (x"97",x"bf",x"7e",x"6e"),
   397 => (x"49",x"c3",x"ff",x"99"),
   398 => (x"c3",x"fe",x"a9",x"05"),
   399 => (x"dd",x"87",x"c0",x"4c"),
   400 => (x"f0",x"e2",x"87",x"d4"),
   401 => (x"66",x"08",x"78",x"d4"),
   402 => (x"66",x"48",x"c4",x"80"),
   403 => (x"d8",x"a6",x"58",x"c1"),
   404 => (x"84",x"c2",x"c0",x"b7"),
   405 => (x"ac",x"04",x"e8",x"87"),
   406 => (x"c1",x"4b",x"4d",x"c1"),
   407 => (x"8b",x"05",x"ff",x"c9"),
   408 => (x"87",x"e3",x"48",x"c3"),
   409 => (x"ff",x"50",x"e7",x"48"),
   410 => (x"c3",x"50",x"75",x"48"),
   411 => (x"26",x"f3",x"f0",x"87"),
   412 => (x"1e",x"73",x"1e",x"71"),
   413 => (x"4b",x"49",x"d8",x"29"),
   414 => (x"c3",x"ff",x"99",x"73"),
   415 => (x"4a",x"c8",x"2a",x"cf"),
   416 => (x"fc",x"c0",x"9a",x"72"),
   417 => (x"b1",x"73",x"4a",x"c8"),
   418 => (x"32",x"c0",x"ff",x"f0"),
   419 => (x"c0",x"c0",x"9a",x"72"),
   420 => (x"b1",x"73",x"4a",x"d8"),
   421 => (x"32",x"ff",x"c0",x"c0"),
   422 => (x"c0",x"c0",x"9a",x"72"),
   423 => (x"b1",x"71",x"48",x"c4"),
   424 => (x"87",x"26",x"4d",x"26"),
   425 => (x"4c",x"26",x"4b",x"26"),
   426 => (x"4f",x"1e",x"73",x"1e"),
   427 => (x"71",x"4b",x"49",x"c8"),
   428 => (x"29",x"c3",x"ff",x"99"),
   429 => (x"73",x"4a",x"c8",x"32"),
   430 => (x"cf",x"fc",x"c0",x"9a"),
   431 => (x"72",x"b1",x"71",x"48"),
   432 => (x"e3",x"87",x"0e",x"5e"),
   433 => (x"5b",x"5c",x"0e",x"71"),
   434 => (x"4b",x"c0",x"4c",x"d0"),
   435 => (x"66",x"48",x"c0",x"b7"),
   436 => (x"a8",x"06",x"c0",x"e3"),
   437 => (x"87",x"13",x"4a",x"cc"),
   438 => (x"66",x"97",x"bf",x"49"),
   439 => (x"cc",x"66",x"48",x"c1"),
   440 => (x"80",x"d0",x"a6",x"58"),
   441 => (x"71",x"b7",x"aa",x"02"),
   442 => (x"c4",x"87",x"c1",x"48"),
   443 => (x"cc",x"87",x"c1",x"84"),
   444 => (x"d0",x"66",x"b7",x"ac"),
   445 => (x"04",x"ff",x"dd",x"87"),
   446 => (x"c0",x"48",x"c2",x"87"),
   447 => (x"26",x"4d",x"26",x"4c"),
   448 => (x"26",x"4b",x"26",x"4f"),
   449 => (x"0e",x"5e",x"5b",x"5c"),
   450 => (x"0e",x"1e",x"c1",x"cc"),
   451 => (x"da",x"48",x"ff",x"78"),
   452 => (x"c1",x"cb",x"ea",x"48"),
   453 => (x"c0",x"78",x"c0",x"e9"),
   454 => (x"de",x"49",x"d9",x"f9"),
   455 => (x"87",x"c1",x"c3",x"e2"),
   456 => (x"1e",x"c0",x"49",x"fb"),
   457 => (x"cf",x"87",x"c4",x"86"),
   458 => (x"70",x"98",x"05",x"c5"),
   459 => (x"87",x"c0",x"48",x"ca"),
   460 => (x"e5",x"87",x"c0",x"4b"),
   461 => (x"c1",x"cc",x"d6",x"48"),
   462 => (x"c1",x"78",x"c8",x"1e"),
   463 => (x"c0",x"e9",x"eb",x"1e"),
   464 => (x"c1",x"c4",x"d8",x"49"),
   465 => (x"fd",x"fb",x"87",x"c8"),
   466 => (x"86",x"70",x"98",x"05"),
   467 => (x"c6",x"87",x"c1",x"cc"),
   468 => (x"d6",x"48",x"c0",x"78"),
   469 => (x"c8",x"1e",x"c0",x"e9"),
   470 => (x"f4",x"1e",x"c1",x"c4"),
   471 => (x"f4",x"49",x"fd",x"e1"),
   472 => (x"87",x"c8",x"86",x"70"),
   473 => (x"98",x"05",x"c6",x"87"),
   474 => (x"c1",x"cc",x"d6",x"48"),
   475 => (x"c0",x"78",x"c8",x"1e"),
   476 => (x"c0",x"e9",x"fd",x"1e"),
   477 => (x"c1",x"c4",x"f4",x"49"),
   478 => (x"fd",x"c7",x"87",x"c8"),
   479 => (x"86",x"70",x"98",x"05"),
   480 => (x"c5",x"87",x"c0",x"48"),
   481 => (x"c9",x"d0",x"87",x"c1"),
   482 => (x"cc",x"d6",x"bf",x"1e"),
   483 => (x"c0",x"ea",x"c6",x"1e"),
   484 => (x"c0",x"e3",x"cb",x"87"),
   485 => (x"c8",x"86",x"c1",x"cc"),
   486 => (x"d6",x"bf",x"02",x"c1"),
   487 => (x"ec",x"87",x"c1",x"c3"),
   488 => (x"e2",x"4a",x"48",x"c6"),
   489 => (x"fe",x"a0",x"4c",x"c1"),
   490 => (x"ca",x"e8",x"bf",x"4b"),
   491 => (x"c1",x"cb",x"e0",x"9f"),
   492 => (x"bf",x"49",x"72",x"7e"),
   493 => (x"c5",x"d6",x"ea",x"a9"),
   494 => (x"05",x"c0",x"cc",x"87"),
   495 => (x"c8",x"a4",x"4a",x"6a"),
   496 => (x"49",x"fa",x"ec",x"87"),
   497 => (x"70",x"4b",x"db",x"87"),
   498 => (x"c7",x"fe",x"a2",x"49"),
   499 => (x"9f",x"69",x"49",x"ca"),
   500 => (x"e9",x"d5",x"a9",x"02"),
   501 => (x"c0",x"cc",x"87",x"c0"),
   502 => (x"e7",x"db",x"49",x"d6"),
   503 => (x"f8",x"87",x"c0",x"48"),
   504 => (x"c7",x"f4",x"87",x"73"),
   505 => (x"1e",x"c0",x"e7",x"f9"),
   506 => (x"1e",x"c0",x"e1",x"f2"),
   507 => (x"87",x"c1",x"c3",x"e2"),
   508 => (x"1e",x"73",x"49",x"f7"),
   509 => (x"ff",x"87",x"cc",x"86"),
   510 => (x"70",x"98",x"05",x"c0"),
   511 => (x"c5",x"87",x"c0",x"48"),
   512 => (x"c7",x"d4",x"87",x"c0"),
   513 => (x"e8",x"d1",x"49",x"d6"),
   514 => (x"cc",x"87",x"c0",x"ea"),
   515 => (x"d9",x"1e",x"c0",x"e1"),
   516 => (x"cd",x"87",x"c8",x"1e"),
   517 => (x"c0",x"ea",x"f1",x"1e"),
   518 => (x"c1",x"c4",x"f4",x"49"),
   519 => (x"fa",x"e3",x"87",x"cc"),
   520 => (x"86",x"70",x"98",x"05"),
   521 => (x"c0",x"c9",x"87",x"c1"),
   522 => (x"cb",x"ea",x"48",x"c1"),
   523 => (x"78",x"c0",x"e4",x"87"),
   524 => (x"c8",x"1e",x"c0",x"ea"),
   525 => (x"fa",x"1e",x"c1",x"c4"),
   526 => (x"d8",x"49",x"fa",x"c5"),
   527 => (x"87",x"c8",x"86",x"70"),
   528 => (x"98",x"02",x"c0",x"cf"),
   529 => (x"87",x"c0",x"e8",x"f8"),
   530 => (x"1e",x"c0",x"e0",x"d2"),
   531 => (x"87",x"c4",x"86",x"c0"),
   532 => (x"48",x"c6",x"c3",x"87"),
   533 => (x"c1",x"cb",x"e0",x"97"),
   534 => (x"bf",x"49",x"c1",x"d5"),
   535 => (x"a9",x"05",x"c0",x"cd"),
   536 => (x"87",x"c1",x"cb",x"e1"),
   537 => (x"97",x"bf",x"49",x"c2"),
   538 => (x"ea",x"a9",x"02",x"c0"),
   539 => (x"c5",x"87",x"c0",x"48"),
   540 => (x"c5",x"e4",x"87",x"c1"),
   541 => (x"c3",x"e2",x"97",x"bf"),
   542 => (x"49",x"c3",x"e9",x"a9"),
   543 => (x"02",x"c0",x"d2",x"87"),
   544 => (x"c1",x"c3",x"e2",x"97"),
   545 => (x"bf",x"49",x"c3",x"eb"),
   546 => (x"a9",x"02",x"c0",x"c5"),
   547 => (x"87",x"c0",x"48",x"c5"),
   548 => (x"c5",x"87",x"c1",x"c3"),
   549 => (x"ed",x"97",x"bf",x"49"),
   550 => (x"99",x"05",x"c0",x"cc"),
   551 => (x"87",x"c1",x"c3",x"ee"),
   552 => (x"97",x"bf",x"49",x"c2"),
   553 => (x"a9",x"02",x"c0",x"c5"),
   554 => (x"87",x"c0",x"48",x"c4"),
   555 => (x"e9",x"87",x"c1",x"c3"),
   556 => (x"ef",x"97",x"bf",x"48"),
   557 => (x"c1",x"cb",x"e6",x"58"),
   558 => (x"c1",x"88",x"c1",x"cb"),
   559 => (x"ea",x"58",x"c1",x"c3"),
   560 => (x"f0",x"97",x"bf",x"49"),
   561 => (x"73",x"81",x"c1",x"c3"),
   562 => (x"f1",x"97",x"bf",x"4a"),
   563 => (x"c8",x"32",x"c1",x"cb"),
   564 => (x"f6",x"48",x"72",x"a1"),
   565 => (x"78",x"c1",x"c3",x"f2"),
   566 => (x"97",x"bf",x"48",x"c1"),
   567 => (x"cc",x"ce",x"58",x"c1"),
   568 => (x"cb",x"ea",x"bf",x"02"),
   569 => (x"c2",x"e0",x"87",x"c8"),
   570 => (x"1e",x"c0",x"e9",x"d5"),
   571 => (x"1e",x"c1",x"c4",x"f4"),
   572 => (x"49",x"f7",x"ce",x"87"),
   573 => (x"c8",x"86",x"70",x"98"),
   574 => (x"02",x"c0",x"c5",x"87"),
   575 => (x"c0",x"48",x"c3",x"d6"),
   576 => (x"87",x"c1",x"cb",x"e2"),
   577 => (x"bf",x"48",x"c4",x"30"),
   578 => (x"c1",x"cc",x"d2",x"58"),
   579 => (x"c1",x"cb",x"e2",x"bf"),
   580 => (x"4a",x"c1",x"cc",x"ca"),
   581 => (x"5a",x"c1",x"c4",x"c7"),
   582 => (x"97",x"bf",x"49",x"c8"),
   583 => (x"31",x"c1",x"c4",x"c6"),
   584 => (x"97",x"bf",x"4b",x"a1"),
   585 => (x"49",x"c1",x"c4",x"c8"),
   586 => (x"97",x"bf",x"4b",x"d0"),
   587 => (x"33",x"73",x"a1",x"49"),
   588 => (x"c1",x"c4",x"c9",x"97"),
   589 => (x"bf",x"4b",x"d8",x"33"),
   590 => (x"73",x"a1",x"49",x"c1"),
   591 => (x"cc",x"d6",x"59",x"c1"),
   592 => (x"cc",x"ca",x"bf",x"91"),
   593 => (x"c1",x"cb",x"f6",x"bf"),
   594 => (x"81",x"c1",x"cb",x"fe"),
   595 => (x"59",x"c1",x"c4",x"cf"),
   596 => (x"97",x"bf",x"4b",x"c8"),
   597 => (x"33",x"c1",x"c4",x"ce"),
   598 => (x"97",x"bf",x"4c",x"a3"),
   599 => (x"4b",x"c1",x"c4",x"d0"),
   600 => (x"97",x"bf",x"4c",x"d0"),
   601 => (x"34",x"74",x"a3",x"4b"),
   602 => (x"c1",x"c4",x"d1",x"97"),
   603 => (x"bf",x"4c",x"cf",x"9c"),
   604 => (x"d8",x"34",x"74",x"a3"),
   605 => (x"4b",x"c1",x"cc",x"c2"),
   606 => (x"5b",x"c2",x"8b",x"73"),
   607 => (x"92",x"c1",x"cc",x"c2"),
   608 => (x"48",x"72",x"a1",x"78"),
   609 => (x"c1",x"ce",x"87",x"c1"),
   610 => (x"c3",x"f4",x"97",x"bf"),
   611 => (x"49",x"c8",x"31",x"c1"),
   612 => (x"c3",x"f3",x"97",x"bf"),
   613 => (x"4a",x"a1",x"49",x"c1"),
   614 => (x"cc",x"d2",x"59",x"c5"),
   615 => (x"31",x"c7",x"ff",x"81"),
   616 => (x"c9",x"29",x"c1",x"cc"),
   617 => (x"ca",x"59",x"c1",x"c3"),
   618 => (x"f9",x"97",x"bf",x"4a"),
   619 => (x"c8",x"32",x"c1",x"c3"),
   620 => (x"f8",x"97",x"bf",x"4b"),
   621 => (x"a2",x"4a",x"c1",x"cc"),
   622 => (x"d6",x"5a",x"c1",x"cc"),
   623 => (x"ca",x"bf",x"92",x"c1"),
   624 => (x"cb",x"f6",x"bf",x"82"),
   625 => (x"c1",x"cc",x"c6",x"5a"),
   626 => (x"c1",x"cb",x"fe",x"48"),
   627 => (x"c0",x"78",x"c1",x"cb"),
   628 => (x"fa",x"48",x"72",x"a1"),
   629 => (x"78",x"c1",x"48",x"26"),
   630 => (x"f4",x"e3",x"87",x"4e"),
   631 => (x"6f",x"20",x"70",x"61"),
   632 => (x"72",x"74",x"69",x"74"),
   633 => (x"69",x"6f",x"6e",x"20"),
   634 => (x"73",x"69",x"67",x"6e"),
   635 => (x"61",x"74",x"75",x"72"),
   636 => (x"65",x"20",x"66",x"6f"),
   637 => (x"75",x"6e",x"64",x"0a"),
   638 => (x"00",x"52",x"65",x"61"),
   639 => (x"64",x"69",x"6e",x"67"),
   640 => (x"20",x"62",x"6f",x"6f"),
   641 => (x"74",x"20",x"73",x"65"),
   642 => (x"63",x"74",x"6f",x"72"),
   643 => (x"20",x"25",x"64",x"0a"),
   644 => (x"00",x"52",x"65",x"61"),
   645 => (x"64",x"20",x"62",x"6f"),
   646 => (x"6f",x"74",x"20",x"73"),
   647 => (x"65",x"63",x"74",x"6f"),
   648 => (x"72",x"20",x"66",x"72"),
   649 => (x"6f",x"6d",x"20",x"66"),
   650 => (x"69",x"72",x"73",x"74"),
   651 => (x"20",x"70",x"61",x"72"),
   652 => (x"74",x"69",x"74",x"69"),
   653 => (x"6f",x"6e",x"0a",x"00"),
   654 => (x"55",x"6e",x"73",x"75"),
   655 => (x"70",x"70",x"6f",x"72"),
   656 => (x"74",x"65",x"64",x"20"),
   657 => (x"70",x"61",x"72",x"74"),
   658 => (x"69",x"74",x"69",x"6f"),
   659 => (x"6e",x"20",x"74",x"79"),
   660 => (x"70",x"65",x"21",x"0d"),
   661 => (x"00",x"46",x"41",x"54"),
   662 => (x"33",x"32",x"20",x"20"),
   663 => (x"20",x"00",x"52",x"65"),
   664 => (x"61",x"64",x"69",x"6e"),
   665 => (x"67",x"20",x"4d",x"42"),
   666 => (x"52",x"0a",x"00",x"46"),
   667 => (x"41",x"54",x"31",x"36"),
   668 => (x"20",x"20",x"20",x"00"),
   669 => (x"46",x"41",x"54",x"33"),
   670 => (x"32",x"20",x"20",x"20"),
   671 => (x"00",x"46",x"41",x"54"),
   672 => (x"31",x"32",x"20",x"20"),
   673 => (x"20",x"00",x"50",x"61"),
   674 => (x"72",x"74",x"69",x"74"),
   675 => (x"69",x"6f",x"6e",x"63"),
   676 => (x"6f",x"75",x"6e",x"74"),
   677 => (x"20",x"25",x"64",x"0a"),
   678 => (x"00",x"48",x"75",x"6e"),
   679 => (x"74",x"69",x"6e",x"67"),
   680 => (x"20",x"66",x"6f",x"72"),
   681 => (x"20",x"66",x"69",x"6c"),
   682 => (x"65",x"73",x"79",x"73"),
   683 => (x"74",x"65",x"6d",x"0a"),
   684 => (x"00",x"46",x"41",x"54"),
   685 => (x"33",x"32",x"20",x"20"),
   686 => (x"20",x"00",x"46",x"41"),
   687 => (x"54",x"31",x"36",x"20"),
   688 => (x"20",x"20",x"00",x"52"),
   689 => (x"65",x"61",x"64",x"69"),
   690 => (x"6e",x"67",x"20",x"64"),
   691 => (x"69",x"72",x"65",x"63"),
   692 => (x"74",x"6f",x"72",x"79"),
   693 => (x"20",x"73",x"65",x"63"),
   694 => (x"74",x"6f",x"72",x"20"),
   695 => (x"25",x"64",x"0a",x"00"),
   696 => (x"66",x"69",x"6c",x"65"),
   697 => (x"20",x"22",x"25",x"73"),
   698 => (x"22",x"20",x"66",x"6f"),
   699 => (x"75",x"6e",x"64",x"0d"),
   700 => (x"00",x"47",x"65",x"74"),
   701 => (x"46",x"41",x"54",x"4c"),
   702 => (x"69",x"6e",x"6b",x"20"),
   703 => (x"72",x"65",x"74",x"75"),
   704 => (x"72",x"6e",x"65",x"64"),
   705 => (x"20",x"25",x"64",x"0a"),
   706 => (x"00",x"43",x"61",x"6e"),
   707 => (x"27",x"74",x"20",x"6f"),
   708 => (x"70",x"65",x"6e",x"20"),
   709 => (x"25",x"73",x"0a",x"00"),
   710 => (x"0e",x"5e",x"5b",x"5c"),
   711 => (x"5d",x"0e",x"71",x"4a"),
   712 => (x"c1",x"cb",x"ea",x"bf"),
   713 => (x"02",x"cc",x"87",x"72"),
   714 => (x"4b",x"c7",x"b7",x"2b"),
   715 => (x"72",x"4c",x"c1",x"ff"),
   716 => (x"9c",x"ca",x"87",x"72"),
   717 => (x"4b",x"c8",x"b7",x"2b"),
   718 => (x"72",x"4c",x"c3",x"ff"),
   719 => (x"9c",x"c1",x"cc",x"da"),
   720 => (x"bf",x"ab",x"02",x"de"),
   721 => (x"87",x"c1",x"c3",x"e2"),
   722 => (x"1e",x"c1",x"cb",x"f6"),
   723 => (x"bf",x"49",x"73",x"81"),
   724 => (x"ea",x"e2",x"87",x"c4"),
   725 => (x"86",x"70",x"98",x"05"),
   726 => (x"c5",x"87",x"c0",x"48"),
   727 => (x"c0",x"f5",x"87",x"c1"),
   728 => (x"cc",x"de",x"5b",x"c1"),
   729 => (x"cb",x"ea",x"bf",x"02"),
   730 => (x"d8",x"87",x"74",x"4a"),
   731 => (x"c4",x"92",x"c1",x"c3"),
   732 => (x"e2",x"82",x"6a",x"49"),
   733 => (x"eb",x"f9",x"87",x"70"),
   734 => (x"49",x"4d",x"cf",x"ff"),
   735 => (x"ff",x"ff",x"ff",x"9d"),
   736 => (x"d0",x"87",x"74",x"4a"),
   737 => (x"c2",x"92",x"c1",x"c3"),
   738 => (x"e2",x"82",x"9f",x"6a"),
   739 => (x"49",x"ec",x"d9",x"87"),
   740 => (x"70",x"4d",x"75",x"48"),
   741 => (x"ed",x"e5",x"87",x"0e"),
   742 => (x"5e",x"5b",x"5c",x"5d"),
   743 => (x"0e",x"f4",x"86",x"71"),
   744 => (x"4c",x"c0",x"4b",x"c1"),
   745 => (x"cc",x"da",x"48",x"ff"),
   746 => (x"78",x"c1",x"cb",x"fe"),
   747 => (x"bf",x"4d",x"c1",x"cc"),
   748 => (x"c2",x"bf",x"7e",x"c1"),
   749 => (x"cb",x"ea",x"bf",x"02"),
   750 => (x"c9",x"87",x"c1",x"cb"),
   751 => (x"e2",x"bf",x"4a",x"c4"),
   752 => (x"32",x"c7",x"87",x"c1"),
   753 => (x"cc",x"c6",x"bf",x"4a"),
   754 => (x"c4",x"32",x"c8",x"a6"),
   755 => (x"5a",x"c8",x"a6",x"48"),
   756 => (x"c0",x"78",x"c4",x"66"),
   757 => (x"48",x"c0",x"a8",x"06"),
   758 => (x"c3",x"cc",x"87",x"c8"),
   759 => (x"66",x"49",x"cf",x"99"),
   760 => (x"05",x"c0",x"e2",x"87"),
   761 => (x"6e",x"1e",x"c0",x"eb"),
   762 => (x"c3",x"1e",x"d1",x"f2"),
   763 => (x"87",x"c1",x"c3",x"e2"),
   764 => (x"1e",x"cc",x"66",x"49"),
   765 => (x"48",x"c1",x"80",x"d0"),
   766 => (x"a6",x"58",x"71",x"e7"),
   767 => (x"f7",x"87",x"cc",x"86"),
   768 => (x"c1",x"c3",x"e2",x"4b"),
   769 => (x"c3",x"87",x"c0",x"e0"),
   770 => (x"83",x"97",x"6b",x"49"),
   771 => (x"99",x"02",x"c2",x"c4"),
   772 => (x"87",x"97",x"6b",x"49"),
   773 => (x"c3",x"e5",x"a9",x"02"),
   774 => (x"c1",x"fa",x"87",x"cb"),
   775 => (x"a3",x"49",x"97",x"69"),
   776 => (x"49",x"d8",x"99",x"05"),
   777 => (x"c1",x"ee",x"87",x"cb"),
   778 => (x"1e",x"c0",x"e0",x"66"),
   779 => (x"1e",x"73",x"49",x"ea"),
   780 => (x"d0",x"87",x"c8",x"86"),
   781 => (x"70",x"98",x"05",x"c1"),
   782 => (x"db",x"87",x"dc",x"a3"),
   783 => (x"4a",x"6a",x"49",x"e8"),
   784 => (x"ee",x"87",x"70",x"4a"),
   785 => (x"c4",x"a4",x"49",x"72"),
   786 => (x"79",x"da",x"a3",x"4a"),
   787 => (x"9f",x"6a",x"49",x"e9"),
   788 => (x"d7",x"87",x"70",x"7e"),
   789 => (x"c1",x"cb",x"ea",x"bf"),
   790 => (x"02",x"d8",x"87",x"d4"),
   791 => (x"a3",x"4a",x"9f",x"6a"),
   792 => (x"49",x"e9",x"c5",x"87"),
   793 => (x"70",x"49",x"c0",x"ff"),
   794 => (x"ff",x"99",x"71",x"48"),
   795 => (x"d0",x"30",x"c8",x"a6"),
   796 => (x"58",x"c5",x"87",x"c4"),
   797 => (x"a6",x"48",x"c0",x"78"),
   798 => (x"c4",x"66",x"4a",x"6e"),
   799 => (x"82",x"c8",x"a4",x"49"),
   800 => (x"72",x"79",x"c0",x"7c"),
   801 => (x"dc",x"66",x"1e",x"c0"),
   802 => (x"eb",x"e0",x"1e",x"cf"),
   803 => (x"d1",x"87",x"c8",x"86"),
   804 => (x"c1",x"48",x"c1",x"ce"),
   805 => (x"87",x"c8",x"66",x"48"),
   806 => (x"c1",x"80",x"cc",x"a6"),
   807 => (x"58",x"c8",x"66",x"48"),
   808 => (x"c4",x"66",x"a8",x"04"),
   809 => (x"fc",x"f4",x"87",x"c1"),
   810 => (x"cb",x"ea",x"bf",x"02"),
   811 => (x"c0",x"f2",x"87",x"75"),
   812 => (x"49",x"f9",x"e4",x"87"),
   813 => (x"70",x"4d",x"1e",x"c0"),
   814 => (x"eb",x"f1",x"1e",x"ce"),
   815 => (x"e1",x"87",x"c8",x"86"),
   816 => (x"75",x"49",x"cf",x"ff"),
   817 => (x"ff",x"ff",x"f8",x"99"),
   818 => (x"a9",x"02",x"d5",x"87"),
   819 => (x"75",x"49",x"c2",x"89"),
   820 => (x"c1",x"cb",x"e2",x"bf"),
   821 => (x"91",x"c1",x"cb",x"fa"),
   822 => (x"bf",x"48",x"71",x"80"),
   823 => (x"70",x"7e",x"fb",x"ec"),
   824 => (x"87",x"c0",x"48",x"f4"),
   825 => (x"8e",x"e8",x"d4",x"87"),
   826 => (x"0e",x"5e",x"5b",x"5c"),
   827 => (x"5d",x"0e",x"1e",x"71"),
   828 => (x"4b",x"1e",x"c1",x"cc"),
   829 => (x"de",x"49",x"fa",x"de"),
   830 => (x"87",x"c4",x"86",x"70"),
   831 => (x"98",x"02",x"c1",x"f5"),
   832 => (x"87",x"c1",x"cc",x"e2"),
   833 => (x"bf",x"49",x"c7",x"ff"),
   834 => (x"81",x"c9",x"29",x"71"),
   835 => (x"7e",x"c0",x"4d",x"4c"),
   836 => (x"6e",x"48",x"c0",x"b7"),
   837 => (x"a8",x"06",x"c1",x"ec"),
   838 => (x"87",x"c1",x"cb",x"fa"),
   839 => (x"bf",x"49",x"c1",x"cc"),
   840 => (x"e6",x"bf",x"4a",x"c2"),
   841 => (x"8a",x"c1",x"cb",x"e2"),
   842 => (x"bf",x"92",x"72",x"a1"),
   843 => (x"49",x"c1",x"cb",x"e6"),
   844 => (x"bf",x"4a",x"74",x"9a"),
   845 => (x"72",x"a1",x"49",x"d4"),
   846 => (x"66",x"1e",x"71",x"e2"),
   847 => (x"f7",x"87",x"c4",x"86"),
   848 => (x"70",x"98",x"05",x"c5"),
   849 => (x"87",x"c0",x"48",x"c1"),
   850 => (x"c0",x"87",x"c1",x"84"),
   851 => (x"c1",x"cb",x"e6",x"bf"),
   852 => (x"49",x"74",x"99",x"05"),
   853 => (x"cc",x"87",x"c1",x"cc"),
   854 => (x"e6",x"bf",x"49",x"f6"),
   855 => (x"fa",x"87",x"c1",x"cc"),
   856 => (x"ea",x"58",x"d4",x"66"),
   857 => (x"48",x"c8",x"c0",x"80"),
   858 => (x"d8",x"a6",x"58",x"c1"),
   859 => (x"85",x"6e",x"b7",x"ad"),
   860 => (x"04",x"fe",x"e5",x"87"),
   861 => (x"cf",x"87",x"73",x"1e"),
   862 => (x"c0",x"ec",x"c9",x"1e"),
   863 => (x"cb",x"e0",x"87",x"c8"),
   864 => (x"86",x"c0",x"48",x"c5"),
   865 => (x"87",x"c1",x"cc",x"e2"),
   866 => (x"bf",x"48",x"26",x"e5"),
   867 => (x"ee",x"87",x"1e",x"f3"),
   868 => (x"48",x"71",x"50",x"48"),
   869 => (x"26",x"4f",x"0e",x"5e"),
   870 => (x"5b",x"5c",x"0e",x"71"),
   871 => (x"4b",x"c0",x"4c",x"13"),
   872 => (x"4a",x"9a",x"02",x"cc"),
   873 => (x"87",x"72",x"49",x"e5"),
   874 => (x"87",x"c1",x"84",x"13"),
   875 => (x"4a",x"9a",x"05",x"f4"),
   876 => (x"87",x"74",x"48",x"c2"),
   877 => (x"87",x"26",x"4d",x"26"),
   878 => (x"4c",x"26",x"4b",x"26"),
   879 => (x"4f",x"0e",x"5e",x"5b"),
   880 => (x"5c",x"5d",x"0e",x"fc"),
   881 => (x"86",x"71",x"4a",x"c0"),
   882 => (x"e0",x"66",x"4c",x"c1"),
   883 => (x"cc",x"ea",x"4b",x"c0"),
   884 => (x"7e",x"72",x"9a",x"05"),
   885 => (x"ce",x"87",x"c1",x"cc"),
   886 => (x"eb",x"4b",x"c1",x"cc"),
   887 => (x"ea",x"48",x"c0",x"f0"),
   888 => (x"50",x"c1",x"ca",x"87"),
   889 => (x"72",x"9a",x"02",x"c0"),
   890 => (x"e5",x"87",x"d4",x"66"),
   891 => (x"4d",x"72",x"1e",x"72"),
   892 => (x"49",x"75",x"4a",x"c9"),
   893 => (x"fd",x"87",x"26",x"4a"),
   894 => (x"c0",x"f9",x"de",x"81"),
   895 => (x"11",x"53",x"72",x"49"),
   896 => (x"75",x"4a",x"c9",x"ee"),
   897 => (x"87",x"70",x"4a",x"c1"),
   898 => (x"8c",x"72",x"9a",x"05"),
   899 => (x"ff",x"de",x"87",x"c0"),
   900 => (x"b7",x"ac",x"06",x"d9"),
   901 => (x"87",x"c0",x"e4",x"66"),
   902 => (x"02",x"c5",x"87",x"c0"),
   903 => (x"f0",x"4a",x"c3",x"87"),
   904 => (x"c0",x"e0",x"4a",x"72"),
   905 => (x"53",x"c1",x"8c",x"c0"),
   906 => (x"b7",x"ac",x"01",x"ff"),
   907 => (x"e7",x"87",x"c1",x"cc"),
   908 => (x"ea",x"ab",x"02",x"dd"),
   909 => (x"87",x"d8",x"66",x"4c"),
   910 => (x"dc",x"66",x"1e",x"c1"),
   911 => (x"8b",x"97",x"6b",x"49"),
   912 => (x"74",x"0f",x"c4",x"86"),
   913 => (x"6e",x"48",x"c1",x"80"),
   914 => (x"70",x"7e",x"c1",x"cc"),
   915 => (x"ea",x"ab",x"05",x"ff"),
   916 => (x"e6",x"87",x"6e",x"48"),
   917 => (x"fc",x"8e",x"26",x"4d"),
   918 => (x"26",x"4c",x"26",x"4b"),
   919 => (x"26",x"4f",x"30",x"31"),
   920 => (x"32",x"33",x"34",x"35"),
   921 => (x"36",x"37",x"38",x"39"),
   922 => (x"41",x"42",x"43",x"44"),
   923 => (x"45",x"46",x"00",x"0e"),
   924 => (x"5e",x"5b",x"5c",x"5d"),
   925 => (x"0e",x"71",x"4b",x"ff"),
   926 => (x"4d",x"13",x"4c",x"9c"),
   927 => (x"02",x"d7",x"87",x"c1"),
   928 => (x"85",x"d4",x"66",x"1e"),
   929 => (x"74",x"49",x"d4",x"66"),
   930 => (x"0f",x"c4",x"86",x"74"),
   931 => (x"a8",x"05",x"c6",x"87"),
   932 => (x"13",x"4c",x"9c",x"05"),
   933 => (x"e9",x"87",x"75",x"48"),
   934 => (x"26",x"4d",x"26",x"4c"),
   935 => (x"26",x"4b",x"26",x"4f"),
   936 => (x"0e",x"5e",x"5b",x"5c"),
   937 => (x"5d",x"0e",x"e8",x"86"),
   938 => (x"71",x"7e",x"c0",x"e8"),
   939 => (x"66",x"4d",x"c0",x"4c"),
   940 => (x"c8",x"a6",x"48",x"c0"),
   941 => (x"78",x"6e",x"97",x"bf"),
   942 => (x"4b",x"6e",x"48",x"c1"),
   943 => (x"80",x"70",x"7e",x"73"),
   944 => (x"9b",x"02",x"c6",x"ce"),
   945 => (x"87",x"c8",x"66",x"02"),
   946 => (x"c5",x"d7",x"87",x"cc"),
   947 => (x"a6",x"48",x"c0",x"78"),
   948 => (x"fc",x"80",x"c0",x"78"),
   949 => (x"73",x"4a",x"c0",x"e0"),
   950 => (x"8a",x"02",x"c3",x"c2"),
   951 => (x"87",x"c3",x"8a",x"02"),
   952 => (x"c2",x"fc",x"87",x"c2"),
   953 => (x"8a",x"02",x"c2",x"e4"),
   954 => (x"87",x"8a",x"02",x"c2"),
   955 => (x"f1",x"87",x"c4",x"8a"),
   956 => (x"02",x"c2",x"eb",x"87"),
   957 => (x"c2",x"8a",x"02",x"c2"),
   958 => (x"e5",x"87",x"c3",x"8a"),
   959 => (x"02",x"c2",x"e7",x"87"),
   960 => (x"d4",x"8a",x"02",x"c0"),
   961 => (x"f4",x"87",x"8a",x"02"),
   962 => (x"c0",x"ff",x"87",x"ca"),
   963 => (x"8a",x"02",x"c0",x"f1"),
   964 => (x"87",x"c1",x"8a",x"02"),
   965 => (x"c1",x"df",x"87",x"8a"),
   966 => (x"02",x"df",x"87",x"c8"),
   967 => (x"8a",x"02",x"c1",x"cd"),
   968 => (x"87",x"c4",x"8a",x"02"),
   969 => (x"c0",x"e3",x"87",x"c3"),
   970 => (x"8a",x"02",x"c0",x"e5"),
   971 => (x"87",x"c2",x"8a",x"02"),
   972 => (x"c8",x"87",x"c3",x"8a"),
   973 => (x"02",x"d3",x"87",x"c1"),
   974 => (x"f9",x"87",x"cc",x"a6"),
   975 => (x"48",x"ca",x"78",x"c2"),
   976 => (x"d2",x"87",x"cc",x"a6"),
   977 => (x"48",x"c2",x"78",x"c2"),
   978 => (x"ca",x"87",x"cc",x"a6"),
   979 => (x"48",x"d0",x"78",x"c2"),
   980 => (x"c2",x"87",x"c0",x"f0"),
   981 => (x"66",x"1e",x"c0",x"f0"),
   982 => (x"66",x"1e",x"c4",x"85"),
   983 => (x"75",x"4a",x"c4",x"8a"),
   984 => (x"6a",x"49",x"fc",x"ca"),
   985 => (x"87",x"c8",x"86",x"70"),
   986 => (x"49",x"a4",x"4c",x"c1"),
   987 => (x"e6",x"87",x"c8",x"a6"),
   988 => (x"48",x"c1",x"78",x"c1"),
   989 => (x"de",x"87",x"c0",x"f0"),
   990 => (x"66",x"1e",x"c4",x"85"),
   991 => (x"75",x"4a",x"c4",x"8a"),
   992 => (x"6a",x"49",x"c0",x"f0"),
   993 => (x"66",x"0f",x"c4",x"86"),
   994 => (x"c1",x"84",x"c1",x"c7"),
   995 => (x"87",x"c0",x"f0",x"66"),
   996 => (x"1e",x"c0",x"e5",x"49"),
   997 => (x"c0",x"f0",x"66",x"0f"),
   998 => (x"c4",x"86",x"c1",x"84"),
   999 => (x"c0",x"f5",x"87",x"c8"),
  1000 => (x"a6",x"48",x"c1",x"78"),
  1001 => (x"c0",x"ed",x"87",x"d0"),
  1002 => (x"a6",x"48",x"c1",x"78"),
  1003 => (x"f8",x"80",x"c1",x"78"),
  1004 => (x"c0",x"e1",x"87",x"c0"),
  1005 => (x"f0",x"ab",x"06",x"db"),
  1006 => (x"87",x"c0",x"f9",x"ab"),
  1007 => (x"03",x"d5",x"87",x"d4"),
  1008 => (x"66",x"49",x"ca",x"91"),
  1009 => (x"73",x"4a",x"c0",x"f0"),
  1010 => (x"8a",x"d4",x"a6",x"48"),
  1011 => (x"72",x"a1",x"78",x"c8"),
  1012 => (x"a6",x"48",x"c1",x"78"),
  1013 => (x"cc",x"66",x"02",x"c1"),
  1014 => (x"e9",x"87",x"c4",x"85"),
  1015 => (x"75",x"49",x"c4",x"89"),
  1016 => (x"a6",x"48",x"69",x"78"),
  1017 => (x"c1",x"e4",x"ab",x"05"),
  1018 => (x"d8",x"87",x"c4",x"66"),
  1019 => (x"48",x"c0",x"b7",x"a8"),
  1020 => (x"03",x"cf",x"87",x"c0"),
  1021 => (x"ed",x"49",x"f6",x"d5"),
  1022 => (x"87",x"c4",x"66",x"48"),
  1023 => (x"c0",x"08",x"88",x"c8"),
  1024 => (x"a6",x"58",x"d0",x"66"),
  1025 => (x"1e",x"d8",x"66",x"1e"),
  1026 => (x"c0",x"f8",x"66",x"1e"),
  1027 => (x"c0",x"f8",x"66",x"1e"),
  1028 => (x"dc",x"66",x"1e",x"d8"),
  1029 => (x"66",x"49",x"f6",x"e4"),
  1030 => (x"87",x"d4",x"86",x"70"),
  1031 => (x"49",x"a4",x"4c",x"c0"),
  1032 => (x"e1",x"87",x"c0",x"e5"),
  1033 => (x"ab",x"05",x"cf",x"87"),
  1034 => (x"d0",x"a6",x"48",x"c0"),
  1035 => (x"78",x"c4",x"80",x"c0"),
  1036 => (x"78",x"f4",x"80",x"c1"),
  1037 => (x"78",x"cc",x"87",x"c0"),
  1038 => (x"f0",x"66",x"1e",x"73"),
  1039 => (x"49",x"c0",x"f0",x"66"),
  1040 => (x"0f",x"c4",x"86",x"6e"),
  1041 => (x"97",x"bf",x"4b",x"6e"),
  1042 => (x"48",x"c1",x"80",x"70"),
  1043 => (x"7e",x"73",x"9b",x"05"),
  1044 => (x"f9",x"f2",x"87",x"74"),
  1045 => (x"48",x"e8",x"8e",x"26"),
  1046 => (x"4d",x"26",x"4c",x"26"),
  1047 => (x"4b",x"26",x"4f",x"1e"),
  1048 => (x"c0",x"1e",x"c0",x"f6"),
  1049 => (x"ce",x"1e",x"d0",x"a6"),
  1050 => (x"1e",x"d0",x"66",x"49"),
  1051 => (x"f8",x"f1",x"87",x"f4"),
  1052 => (x"8e",x"26",x"4f",x"1e"),
  1053 => (x"73",x"1e",x"72",x"9a"),
  1054 => (x"02",x"c0",x"e7",x"87"),
  1055 => (x"c0",x"48",x"c1",x"4b"),
  1056 => (x"72",x"a9",x"06",x"d1"),
  1057 => (x"87",x"72",x"82",x"06"),
  1058 => (x"c9",x"87",x"73",x"83"),
  1059 => (x"72",x"a9",x"01",x"f4"),
  1060 => (x"87",x"c3",x"87",x"c1"),
  1061 => (x"b2",x"3a",x"72",x"a9"),
  1062 => (x"03",x"89",x"73",x"80"),
  1063 => (x"07",x"c1",x"2a",x"2b"),
  1064 => (x"05",x"f3",x"87",x"26"),
  1065 => (x"4b",x"26",x"4f",x"1e"),
  1066 => (x"75",x"1e",x"c4",x"4d"),
  1067 => (x"71",x"b7",x"a1",x"04"),
  1068 => (x"ff",x"b9",x"c1",x"81"),
  1069 => (x"c3",x"bd",x"07",x"72"),
  1070 => (x"b7",x"a2",x"04",x"ff"),
  1071 => (x"ba",x"c1",x"82",x"c1"),
  1072 => (x"bd",x"07",x"fe",x"ee"),
  1073 => (x"87",x"c1",x"2d",x"04"),
  1074 => (x"ff",x"b8",x"c1",x"80"),
  1075 => (x"07",x"2d",x"04",x"ff"),
  1076 => (x"b9",x"c1",x"81",x"07"),
  1077 => (x"26",x"4d",x"26",x"4f"),
	others => (others => x"00")
);

-- Xilinx XST attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "no_rw_check";

-- Altera Quartus attributes
attribute ramstyle: string;
attribute ramstyle of ram: signal is "no_rw_check";

signal q_local : word_t;
signal q2_local : word_t;

begin
    
	process(clk,q_local)
	begin

		q(31 downto 24)<=q_local(0);
		q(23 downto 16)<=q_local(1);
		q(15 downto 8)<=q_local(2);
		q(7 downto 0)<=q_local(3);

		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel(3) = '1') then
					ram(to_integer(unsigned(addr)))(3) <= d(7 downto 0);
				end if;
				if bytesel(2) = '1' then
					ram(to_integer(unsigned(addr)))(2) <= d(15 downto 8);
				end if;
				if bytesel(1) = '1' then
					ram(to_integer(unsigned(addr)))(1) <= d(23 downto 16);
				end if;
				if bytesel(0) = '1' then
					ram(to_integer(unsigned(addr)))(0) <= d(31 downto 24);
				end if;
			end if;
			q_local <= ram(to_integer(unsigned(addr)));
		end if;
	end process;

	-- Second port
	
	process(clk,q2_local)
	begin

		q2(31 downto 24)<=q2_local(0);
		q2(23 downto 16)<=q2_local(1);
		q2(15 downto 8)<=q2_local(2);
		q2(7 downto 0)<=q2_local(3);

		if(rising_edge(clk)) then 
			if(we2 = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel2(3) = '1') then
					ram(to_integer(unsigned(addr2)))(3) <= d2(7 downto 0);
				end if;
				if bytesel2(2) = '1' then
					ram(to_integer(unsigned(addr2)))(2) <= d2(15 downto 8);
				end if;
				if bytesel2(1) = '1' then
					ram(to_integer(unsigned(addr2)))(1) <= d2(23 downto 16);
				end if;
				if bytesel2(0) = '1' then
					ram(to_integer(unsigned(addr2)))(0) <= d2(31 downto 24);
				end if;
			end if;
			q2_local <= ram(to_integer(unsigned(addr2)));
		end if;
	end process;

end arch;

